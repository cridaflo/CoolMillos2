// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition"

// DATE "12/06/2018 09:08:56"

// 
// Device: Altera EP4CE22F17C6 Package FBGA256
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module niosII (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	adc_0_sclk,
	adc_0_cs_n,
	adc_0_dout,
	adc_0_din,
	clk_clk,
	epcs_dclk,
	epcs_sce,
	epcs_sdo,
	epcs_data0,
	port_gpio_0_export,
	port_key_export,
	port_led_export,
	port_sw_export,
	ram_clk_clk,
	reset_reset_n,
	rs232_0_RXD,
	rs232_0_TXD,
	rs232_1_RXD,
	rs232_1_TXD,
	sdram_addr,
	sdram_ba,
	sdram_cas_n,
	sdram_cke,
	sdram_cs_n,
	sdram_dq,
	sdram_dqm,
	sdram_ras_n,
	sdram_we_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
output 	adc_0_sclk;
output 	adc_0_cs_n;
input 	adc_0_dout;
output 	adc_0_din;
input 	clk_clk;
output 	epcs_dclk;
output 	epcs_sce;
output 	epcs_sdo;
input 	epcs_data0;
inout 	[31:0] port_gpio_0_export;
input 	[1:0] port_key_export;
output 	[7:0] port_led_export;
input 	[3:0] port_sw_export;
output 	ram_clk_clk;
input 	reset_reset_n;
input 	rs232_0_RXD;
output 	rs232_0_TXD;
input 	rs232_1_RXD;
output 	rs232_1_TXD;
output 	[12:0] sdram_addr;
output 	[1:0] sdram_ba;
output 	sdram_cas_n;
output 	sdram_cke;
output 	sdram_cs_n;
inout 	[15:0] sdram_dq;
output 	[1:0] sdram_dqm;
output 	sdram_ras_n;
output 	sdram_we_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sys_pll|sd1|wire_pll7_clk[0] ;
wire \sys_pll|sd1|wire_pll7_clk[1] ;
wire \sdram|m_addr[0]~q ;
wire \sdram|m_addr[1]~q ;
wire \sdram|m_addr[2]~q ;
wire \sdram|m_addr[3]~q ;
wire \sdram|m_addr[4]~q ;
wire \sdram|m_addr[5]~q ;
wire \sdram|m_addr[6]~q ;
wire \sdram|m_addr[7]~q ;
wire \sdram|m_addr[8]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|sr[0]~q ;
wire \cpu|cpu|W_alu_result[6]~q ;
wire \cpu|cpu|W_alu_result[26]~q ;
wire \cpu|cpu|W_alu_result[25]~q ;
wire \cpu|cpu|W_alu_result[24]~q ;
wire \cpu|cpu|W_alu_result[23]~q ;
wire \cpu|cpu|W_alu_result[22]~q ;
wire \cpu|cpu|W_alu_result[21]~q ;
wire \cpu|cpu|W_alu_result[20]~q ;
wire \cpu|cpu|W_alu_result[19]~q ;
wire \cpu|cpu|W_alu_result[18]~q ;
wire \cpu|cpu|W_alu_result[17]~q ;
wire \cpu|cpu|W_alu_result[16]~q ;
wire \cpu|cpu|W_alu_result[15]~q ;
wire \cpu|cpu|W_alu_result[14]~q ;
wire \cpu|cpu|W_alu_result[13]~q ;
wire \cpu|cpu|W_alu_result[12]~q ;
wire \cpu|cpu|W_alu_result[11]~q ;
wire \cpu|cpu|W_alu_result[10]~q ;
wire \cpu|cpu|W_alu_result[5]~q ;
wire \cpu|cpu|W_alu_result[7]~q ;
wire \cpu|cpu|W_alu_result[9]~q ;
wire \cpu|cpu|W_alu_result[8]~q ;
wire \cpu|cpu|W_alu_result[4]~q ;
wire \cpu|cpu|W_alu_result[3]~q ;
wire \cpu|cpu|W_alu_result[2]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|byteen_reg[0]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|byteen_reg[1]~q ;
wire \sdram|oe~q ;
wire \cpu|cpu|d_writedata[24]~q ;
wire \cpu|cpu|d_writedata[25]~q ;
wire \cpu|cpu|d_writedata[26]~q ;
wire \cpu|cpu|d_writedata[27]~q ;
wire \cpu|cpu|d_writedata[28]~q ;
wire \cpu|cpu|d_writedata[29]~q ;
wire \cpu|cpu|d_writedata[30]~q ;
wire \cpu|cpu|d_writedata[31]~q ;
wire \rs232_0|readdata[0]~q ;
wire \rs232_1|readdata[0]~q ;
wire \rs232_1|irq~q ;
wire \rs232_0|irq~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[4]~q ;
wire \rs232_0|readdata[1]~q ;
wire \rs232_1|readdata[1]~q ;
wire \rs232_0|readdata[23]~q ;
wire \rs232_1|readdata[23]~q ;
wire \rs232_1|readdata[22]~q ;
wire \rs232_0|readdata[22]~q ;
wire \rs232_1|readdata[21]~q ;
wire \rs232_0|readdata[21]~q ;
wire \rs232_1|readdata[20]~q ;
wire \rs232_0|readdata[20]~q ;
wire \rs232_1|readdata[19]~q ;
wire \rs232_0|readdata[19]~q ;
wire \rs232_1|readdata[18]~q ;
wire \rs232_0|readdata[18]~q ;
wire \rs232_1|readdata[17]~q ;
wire \rs232_0|readdata[17]~q ;
wire \rs232_1|readdata[16]~q ;
wire \rs232_0|readdata[16]~q ;
wire \adc_0|ADC_CTRL|sclk~q ;
wire \adc_0|ADC_CTRL|cs_n~2_combout ;
wire \adc_0|ADC_CTRL|addr_shift_reg[5]~q ;
wire \epcs|the_niosII_epcs_sub|SCLK_reg~q ;
wire \epcs|the_niosII_epcs_sub|SS_n~0_combout ;
wire \epcs|the_niosII_epcs_sub|shift_reg[7]~q ;
wire \port_led|data_out[0]~q ;
wire \port_led|data_out[1]~q ;
wire \port_led|data_out[2]~q ;
wire \port_led|data_out[3]~q ;
wire \port_led|data_out[4]~q ;
wire \port_led|data_out[5]~q ;
wire \port_led|data_out[6]~q ;
wire \port_led|data_out[7]~q ;
wire \rs232_0|RS232_Out_Serializer|serial_data_out~q ;
wire \rs232_1|RS232_Out_Serializer|serial_data_out~q ;
wire \sdram|m_addr[9]~q ;
wire \sdram|m_addr[10]~q ;
wire \sdram|m_addr[11]~q ;
wire \sdram|m_addr[12]~q ;
wire \sdram|m_bank[0]~q ;
wire \sdram|m_bank[1]~q ;
wire \sdram|m_cmd[1]~q ;
wire \sdram|m_cmd[3]~q ;
wire \sdram|m_dqm[0]~q ;
wire \sdram|m_dqm[1]~q ;
wire \sdram|m_cmd[2]~q ;
wire \sdram|m_cmd[0]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|ir_out[0]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|ir_out[1]~q ;
wire \jtag|niosII_jtag_alt_jtag_atlantic|tdo~q ;
wire \rst_controller|r_sync_rst~q ;
wire \rst_controller_001|r_sync_rst~q ;
wire \mm_interconnect_0|cmd_mux_010|saved_grant[0]~q ;
wire \mm_interconnect_0|cmd_mux_010|saved_grant[1]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[38]~q ;
wire \mm_interconnect_0|cmd_mux_010|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_010|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_010|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~0_combout ;
wire \sdram|the_niosII_sdram_input_efifo_module|entries[1]~q ;
wire \sdram|the_niosII_sdram_input_efifo_module|entries[0]~q ;
wire \mm_interconnect_0|adc_0_adc_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \cpu|cpu|d_read~q ;
wire \mm_interconnect_0|cpu_data_master_translator|read_accepted~q ;
wire \mm_interconnect_0|cpu_data_master_agent|hold_waitrequest~q ;
wire \cpu|cpu|d_write~q ;
wire \mm_interconnect_0|cpu_data_master_translator|write_accepted~q ;
wire \mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ;
wire \mm_interconnect_0|router|Equal3~6_combout ;
wire \mm_interconnect_0|adc_0_adc_slave_agent|m0_read~combout ;
wire \mm_interconnect_0|timer_0_s1_agent|m0_write~0_combout ;
wire \timer_0|read_mux_out~0_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~1_combout ;
wire \mm_interconnect_0|epcs_epcs_control_port_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|epcs_epcs_control_port_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|cmd_mux_010|src_valid~0_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_valid~1_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_data[46]~combout ;
wire \mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[65]~q ;
wire \epcs|the_niosII_epcs_sub|p1_wr_strobe~1_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~2_combout ;
wire \cpu|cpu|d_writedata[0]~q ;
wire \port_led|data~0_combout ;
wire \cpu|cpu|d_byteenable[0]~q ;
wire \timer_0|Equal6~0_combout ;
wire \mm_interconnect_0|router|Equal9~0_combout ;
wire \mm_interconnect_0|port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg~0_combout ;
wire \cpu|cpu|d_writedata[1]~q ;
wire \port_led|data~3_combout ;
wire \cpu|cpu|d_writedata[2]~q ;
wire \port_led|data~4_combout ;
wire \cpu|cpu|d_writedata[3]~q ;
wire \port_led|data~5_combout ;
wire \cpu|cpu|d_writedata[4]~q ;
wire \port_led|data~6_combout ;
wire \cpu|cpu|d_writedata[5]~q ;
wire \port_led|data~7_combout ;
wire \cpu|cpu|d_writedata[6]~q ;
wire \port_led|data~8_combout ;
wire \cpu|cpu|d_writedata[7]~q ;
wire \port_led|data~9_combout ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[0]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_toggle_flopped~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \mm_interconnect_0|sys_pll_pll_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \sys_pll|wire_pfdena_reg_ena~0_combout ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[65]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[38]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[39]~q ;
wire \rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \mm_interconnect_0|cmd_mux_012|saved_grant[0]~q ;
wire \cpu|cpu|d_byteenable[1]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|use_reg~q ;
wire \mm_interconnect_0|cmd_mux_012|saved_grant[1]~q ;
wire \mm_interconnect_0|sdram_s1_agent|WideOr0~2_combout ;
wire \sdram|the_niosII_sdram_input_efifo_module|Equal0~0_combout ;
wire \cpu|cpu|i_read~q ;
wire \cpu|cpu|F_pc[24]~q ;
wire \cpu|cpu|F_pc[23]~q ;
wire \cpu|cpu|F_pc[22]~q ;
wire \cpu|cpu|F_pc[21]~q ;
wire \cpu|cpu|F_pc[20]~q ;
wire \cpu|cpu|F_pc[19]~q ;
wire \cpu|cpu|F_pc[18]~q ;
wire \cpu|cpu|F_pc[17]~q ;
wire \cpu|cpu|F_pc[16]~q ;
wire \cpu|cpu|F_pc[15]~q ;
wire \cpu|cpu|F_pc[14]~q ;
wire \cpu|cpu|F_pc[13]~q ;
wire \cpu|cpu|F_pc[12]~q ;
wire \cpu|cpu|F_pc[11]~q ;
wire \cpu|cpu|F_pc[10]~q ;
wire \mm_interconnect_0|router|Equal1~0_combout ;
wire \mm_interconnect_0|router|Equal4~1_combout ;
wire \mm_interconnect_0|cmd_mux_012|WideOr1~combout ;
wire \mm_interconnect_0|sdram_s1_agent|m0_write~2_combout ;
wire \mm_interconnect_0|sdram_s1_agent_rsp_fifo|mem_used[7]~q ;
wire \mm_interconnect_0|cmd_mux_012|src_data[66]~combout ;
wire \cpu|cpu|F_pc[8]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[28]~0_combout ;
wire \mm_interconnect_0|cmd_mux_012|src_valid~0_combout ;
wire \mm_interconnect_0|cmd_demux|src12_valid~0_combout ;
wire \mm_interconnect_0|sdram_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[42]~1_combout ;
wire \cpu|cpu|F_pc[9]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[29]~2_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[31]~3_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[30]~4_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[33]~5_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[32]~6_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[35]~7_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[34]~8_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[37]~9_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[36]~10_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[39]~11_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[38]~12_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[41]~13_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[40]~14_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[19]~15_combout ;
wire \cpu|cpu|F_pc[0]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[20]~16_combout ;
wire \cpu|cpu|F_pc[1]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[21]~17_combout ;
wire \cpu|cpu|F_pc[2]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[22]~18_combout ;
wire \cpu|cpu|F_pc[3]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[23]~19_combout ;
wire \cpu|cpu|F_pc[4]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[24]~20_combout ;
wire \cpu|cpu|F_pc[5]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[25]~21_combout ;
wire \cpu|cpu|F_pc[6]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[26]~22_combout ;
wire \cpu|cpu|F_pc[7]~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[27]~23_combout ;
wire \port_gpio_0|data_out[0]~q ;
wire \port_gpio_0|direction[0]~q ;
wire \port_gpio_0|data_out[1]~q ;
wire \port_gpio_0|direction[1]~q ;
wire \port_gpio_0|data_out[2]~q ;
wire \port_gpio_0|direction[2]~q ;
wire \port_gpio_0|data_out[3]~q ;
wire \port_gpio_0|direction[3]~q ;
wire \port_gpio_0|data_out[4]~q ;
wire \port_gpio_0|direction[4]~q ;
wire \port_gpio_0|data_out[5]~q ;
wire \port_gpio_0|direction[5]~q ;
wire \port_gpio_0|data_out[6]~q ;
wire \port_gpio_0|direction[6]~q ;
wire \port_gpio_0|data_out[7]~q ;
wire \port_gpio_0|direction[7]~q ;
wire \port_gpio_0|data_out[8]~q ;
wire \port_gpio_0|direction[8]~q ;
wire \port_gpio_0|data_out[9]~q ;
wire \port_gpio_0|direction[9]~q ;
wire \port_gpio_0|data_out[10]~q ;
wire \port_gpio_0|direction[10]~q ;
wire \port_gpio_0|data_out[11]~q ;
wire \port_gpio_0|direction[11]~q ;
wire \port_gpio_0|data_out[12]~q ;
wire \port_gpio_0|direction[12]~q ;
wire \port_gpio_0|data_out[13]~q ;
wire \port_gpio_0|direction[13]~q ;
wire \port_gpio_0|data_out[14]~q ;
wire \port_gpio_0|direction[14]~q ;
wire \port_gpio_0|data_out[15]~q ;
wire \port_gpio_0|direction[15]~q ;
wire \port_gpio_0|data_out[16]~q ;
wire \port_gpio_0|direction[16]~q ;
wire \port_gpio_0|data_out[17]~q ;
wire \port_gpio_0|direction[17]~q ;
wire \port_gpio_0|data_out[18]~q ;
wire \port_gpio_0|direction[18]~q ;
wire \port_gpio_0|data_out[19]~q ;
wire \port_gpio_0|direction[19]~q ;
wire \port_gpio_0|data_out[20]~q ;
wire \port_gpio_0|direction[20]~q ;
wire \port_gpio_0|data_out[21]~q ;
wire \port_gpio_0|direction[21]~q ;
wire \port_gpio_0|data_out[22]~q ;
wire \port_gpio_0|direction[22]~q ;
wire \port_gpio_0|data_out[23]~q ;
wire \port_gpio_0|direction[23]~q ;
wire \port_gpio_0|data_out[24]~q ;
wire \port_gpio_0|direction[24]~q ;
wire \port_gpio_0|data_out[25]~q ;
wire \port_gpio_0|direction[25]~q ;
wire \port_gpio_0|data_out[26]~q ;
wire \port_gpio_0|direction[26]~q ;
wire \port_gpio_0|data_out[27]~q ;
wire \port_gpio_0|direction[27]~q ;
wire \port_gpio_0|data_out[28]~q ;
wire \port_gpio_0|direction[28]~q ;
wire \port_gpio_0|data_out[29]~q ;
wire \port_gpio_0|direction[29]~q ;
wire \port_gpio_0|data_out[30]~q ;
wire \port_gpio_0|direction[30]~q ;
wire \port_gpio_0|data_out[31]~q ;
wire \port_gpio_0|direction[31]~q ;
wire \sdram|m_data[0]~q ;
wire \sdram|m_data[1]~q ;
wire \sdram|m_data[2]~q ;
wire \sdram|m_data[3]~q ;
wire \sdram|m_data[4]~q ;
wire \sdram|m_data[5]~q ;
wire \sdram|m_data[6]~q ;
wire \sdram|m_data[7]~q ;
wire \sdram|m_data[8]~q ;
wire \sdram|m_data[9]~q ;
wire \sdram|m_data[10]~q ;
wire \sdram|m_data[11]~q ;
wire \sdram|m_data[12]~q ;
wire \sdram|m_data[13]~q ;
wire \sdram|m_data[14]~q ;
wire \sdram|m_data[15]~q ;
wire \adc_0|always0~1_combout ;
wire \adc_0|waitrequest~0_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][84]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][66]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|port_gpio_0_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|sys_id_control_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rsp_fifo|mem[0][54]~q ;
wire \mm_interconnect_0|rsp_demux_012|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|timer_0_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|timer_0_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|timer_0_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg~2_combout ;
wire \mm_interconnect_0|port_sw_avalon_parallel_port_slave_agent_rsp_fifo|write~2_combout ;
wire \mm_interconnect_0|router|Equal12~1_combout ;
wire \mm_interconnect_0|rs232_0_avalon_rs232_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_009|saved_grant[0]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cpu_data_master_translator|av_waitrequest~1_combout ;
wire \timer_0|Equal6~1_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_data[66]~combout ;
wire \mm_interconnect_0|epcs_epcs_control_port_translator|av_begintransfer~0_combout ;
wire \cpu|cpu|d_writedata[10]~q ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~4_combout ;
wire \jtag|niosII_jtag_alt_jtag_atlantic|rst1~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[66]~q ;
wire \cpu|cpu|d_byteenable[2]~q ;
wire \cpu|cpu|d_byteenable[3]~q ;
wire \mm_interconnect_0|rsp_demux_009|src1_valid~0_combout ;
wire \mm_interconnect_0|cpu_instruction_master_translator|read_accepted~2_combout ;
wire \mm_interconnect_0|rsp_demux_012|src1_valid~0_combout ;
wire \cpu|cpu|hbreak_enabled~q ;
wire \mm_interconnect_0|port_gpio_0_avalon_parallel_port_slave_translator|read_latency_shift_reg~0_combout ;
wire \cpu|cpu|d_writedata[8]~q ;
wire \cpu|cpu|d_writedata[9]~q ;
wire \cpu|cpu|d_writedata[11]~q ;
wire \cpu|cpu|d_writedata[12]~q ;
wire \cpu|cpu|d_writedata[13]~q ;
wire \cpu|cpu|d_writedata[14]~q ;
wire \cpu|cpu|d_writedata[15]~q ;
wire \cpu|cpu|d_writedata[16]~q ;
wire \cpu|cpu|d_writedata[17]~q ;
wire \cpu|cpu|d_writedata[18]~q ;
wire \cpu|cpu|d_writedata[19]~q ;
wire \cpu|cpu|d_writedata[20]~q ;
wire \cpu|cpu|d_writedata[21]~q ;
wire \cpu|cpu|d_writedata[22]~q ;
wire \cpu|cpu|d_writedata[23]~q ;
wire \mm_interconnect_0|cmd_mux_009|WideOr1~combout ;
wire \mm_interconnect_0|port_key_avalon_parallel_port_slave_agent_rsp_fifo|write~0_combout ;
wire \mm_interconnect_0|router|Equal12~2_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent|rf_source_valid~0_combout ;
wire \mm_interconnect_0|cpu_data_master_translator|uav_write~0_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~5_combout ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_valid~combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[0]~q ;
wire \mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[0]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[0]~q ;
wire \mm_interconnect_0|sdram_s1_agent|uncompressor|source_addr[1]~0_combout ;
wire \cpu|cpu|F_iw[0]~5_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[1]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[1]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~16_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[2]~q ;
wire \mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[2]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[2]~q ;
wire \cpu|cpu|F_iw[2]~10_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[3]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[3]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~17_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[4]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[4]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~18_combout ;
wire \rs232_0|data_to_uart[0]~q ;
wire \port_led|data~10_combout ;
wire \mm_interconnect_0|rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg~1_combout ;
wire \rst_controller|r_early_rst~q ;
wire \jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[0]~24_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[1]~25_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[2]~26_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[3]~27_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[4]~28_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[5]~29_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[6]~30_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[7]~31_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[8]~32_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[9]~33_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[10]~34_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[11]~35_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[12]~36_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[13]~37_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[14]~38_combout ;
wire \mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[15]~39_combout ;
wire \timer_0|period_l_wr_strobe~2_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[46]~combout ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_toggle_flopped~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[11]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[11]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[11]~19_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[13]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[13]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[13]~20_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[16]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~0_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[12]~q ;
wire \mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[12]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[12]~q ;
wire \cpu|cpu|F_iw[12]~23_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[5]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[5]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~21_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[14]~q ;
wire \mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[14]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[14]~q ;
wire \cpu|cpu|F_iw[14]~28_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[15]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[15]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[15]~22_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[10]~q ;
wire \mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[10]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[10]~q ;
wire \cpu|cpu|F_iw[10]~33_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[9]~q ;
wire \mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[9]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[9]~q ;
wire \cpu|cpu|F_iw[9]~36_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[8]~q ;
wire \mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[8]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[8]~q ;
wire \cpu|cpu|F_iw[8]~39_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[7]~q ;
wire \mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[7]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[7]~q ;
wire \cpu|cpu|F_iw[7]~42_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[6]~q ;
wire \mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[6]~q ;
wire \mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[6]~q ;
wire \cpu|cpu|F_iw[6]~45_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[21]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[30]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[29]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[28]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[27]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[26]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[25]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[24]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[23]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[22]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[20]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[19]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[18]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[17]~q ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~6_combout ;
wire \port_led|readdata[0]~q ;
wire \port_sw|readdata[0]~q ;
wire \port_key|readdata[0]~q ;
wire \port_gpio_0|readdata[0]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_valid~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~30_combout ;
wire \irq_synchronizer_001|sync|sync[0].u|dreg[1]~q ;
wire \timer_0|timeout_occurred~q ;
wire \timer_0|control_register[0]~q ;
wire \irq_synchronizer|sync|sync[0].u|dreg[1]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[0]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[1]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[2]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[3]~q ;
wire \port_led|readdata[1]~q ;
wire \port_sw|readdata[1]~q ;
wire \port_key|readdata[1]~q ;
wire \port_gpio_0|readdata[1]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~38_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~39_combout ;
wire \port_led|readdata[2]~q ;
wire \port_gpio_0|readdata[2]~q ;
wire \port_sw|readdata[2]~q ;
wire \rs232_1|readdata[2]~q ;
wire \rs232_0|readdata[2]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~45_combout ;
wire \port_led|readdata[3]~q ;
wire \port_gpio_0|readdata[3]~q ;
wire \port_sw|readdata[3]~q ;
wire \rs232_1|readdata[3]~q ;
wire \rs232_0|readdata[3]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~52_combout ;
wire \port_led|readdata[4]~q ;
wire \rs232_0|readdata[4]~q ;
wire \port_gpio_0|readdata[4]~q ;
wire \rs232_1|readdata[4]~q ;
wire \mm_interconnect_0|sys_id_control_slave_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~58_combout ;
wire \port_led|readdata[5]~q ;
wire \rs232_0|readdata[5]~q ;
wire \port_gpio_0|readdata[5]~q ;
wire \rs232_1|readdata[5]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~64_combout ;
wire \port_led|readdata[6]~q ;
wire \rs232_0|readdata[6]~q ;
wire \port_gpio_0|readdata[6]~q ;
wire \rs232_1|readdata[6]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[6]~70_combout ;
wire \port_led|readdata[7]~q ;
wire \rs232_0|readdata[7]~q ;
wire \port_gpio_0|readdata[7]~q ;
wire \rs232_1|readdata[7]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[7]~76_combout ;
wire \rs232_0|data_to_uart[1]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[32]~combout ;
wire \jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \mm_interconnect_0|crosser|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \jtag|av_waitrequest~q ;
wire \mm_interconnect_0|jtag_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[66]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[38]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[7]~q ;
wire \sdram|za_valid~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[11]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[13]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[16]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[12]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[5]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[14]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[15]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[10]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[31]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[9]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[8]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[7]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[6]~q ;
wire \port_gpio_0|readdata[26]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[26]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[21]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[30]~q ;
wire \port_gpio_0|readdata[25]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[25]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~5_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[29]~q ;
wire \port_gpio_0|readdata[24]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[24]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[28]~q ;
wire \port_gpio_0|readdata[23]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~9_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[27]~q ;
wire \port_gpio_0|readdata[22]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~14_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[26]~q ;
wire \port_gpio_0|readdata[21]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~19_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[25]~q ;
wire \port_gpio_0|readdata[20]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~24_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[24]~q ;
wire \port_gpio_0|readdata[19]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~29_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[23]~q ;
wire \port_gpio_0|readdata[18]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~34_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[22]~q ;
wire \port_gpio_0|readdata[17]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~39_combout ;
wire \port_gpio_0|readdata[16]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~44_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[20]~q ;
wire \port_gpio_0|readdata[15]~q ;
wire \rs232_1|readdata[15]~q ;
wire \rs232_0|readdata[15]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[15]~82_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[19]~q ;
wire \port_gpio_0|readdata[14]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[14]~85_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[18]~q ;
wire \port_gpio_0|readdata[13]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[13]~89_combout ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[17]~q ;
wire \port_gpio_0|readdata[12]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[12]~92_combout ;
wire \port_gpio_0|readdata[11]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[11]~96_combout ;
wire \port_gpio_0|readdata[10]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[10]~101_combout ;
wire \port_gpio_0|readdata[9]~q ;
wire \rs232_1|readdata[9]~q ;
wire \rs232_0|readdata[9]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[9]~107_combout ;
wire \port_gpio_0|readdata[8]~q ;
wire \rs232_1|readdata[8]~q ;
wire \rs232_0|readdata[8]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[8]~113_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~7_combout ;
wire \mm_interconnect_0|adc_0_adc_slave_translator|av_readdata_pre[0]~0_combout ;
wire \adc_0|readdata[0]~4_combout ;
wire \timer_0|readdata[0]~q ;
wire \adc_0|readdata[1]~9_combout ;
wire \timer_0|readdata[1]~q ;
wire \adc_0|readdata[2]~14_combout ;
wire \timer_0|readdata[2]~q ;
wire \adc_0|readdata[3]~19_combout ;
wire \timer_0|readdata[3]~q ;
wire \adc_0|readdata[4]~24_combout ;
wire \timer_0|readdata[4]~q ;
wire \adc_0|readdata[5]~29_combout ;
wire \timer_0|readdata[5]~q ;
wire \adc_0|readdata[6]~34_combout ;
wire \timer_0|readdata[6]~q ;
wire \adc_0|readdata[7]~39_combout ;
wire \timer_0|readdata[7]~q ;
wire \rs232_0|data_to_uart[2]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~2_combout ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[65]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[0]~q ;
wire \jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \port_gpio_0|readdata[27]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[27]~q ;
wire \port_gpio_0|readdata[28]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[28]~q ;
wire \port_gpio_0|readdata[29]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[29]~q ;
wire \port_gpio_0|readdata[30]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[30]~q ;
wire \port_gpio_0|readdata[31]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[31]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[31]~q ;
wire \adc_0|readdata[15]~40_combout ;
wire \timer_0|readdata[15]~q ;
wire \timer_0|readdata[14]~q ;
wire \timer_0|readdata[13]~q ;
wire \timer_0|readdata[12]~q ;
wire \adc_0|readdata[11]~45_combout ;
wire \timer_0|readdata[11]~q ;
wire \timer_0|readdata[10]~q ;
wire \adc_0|readdata[10]~50_combout ;
wire \adc_0|readdata[9]~55_combout ;
wire \timer_0|readdata[9]~q ;
wire \adc_0|readdata[8]~60_combout ;
wire \timer_0|readdata[8]~q ;
wire \cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_oci_debug|resetrequest~q ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~8_combout ;
wire \rs232_0|RS232_In_Deserializer|comb~1_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~5_combout ;
wire \epcs|readdata[0]~0_combout ;
wire \sdram|za_data[0]~q ;
wire \epcs|readdata[1]~1_combout ;
wire \sdram|za_data[1]~q ;
wire \epcs|readdata[2]~2_combout ;
wire \sdram|za_data[2]~q ;
wire \epcs|readdata[3]~3_combout ;
wire \sdram|za_data[3]~q ;
wire \epcs|readdata[4]~4_combout ;
wire \sdram|za_data[4]~q ;
wire \rs232_0|data_to_uart[3]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[1]~q ;
wire \epcs|readdata[11]~5_combout ;
wire \sdram|za_data[11]~q ;
wire \epcs|readdata[13]~6_combout ;
wire \sdram|za_data[13]~q ;
wire \epcs|readdata[16]~7_combout ;
wire \epcs|readdata[12]~8_combout ;
wire \sdram|za_data[12]~q ;
wire \epcs|readdata[5]~9_combout ;
wire \sdram|za_data[5]~q ;
wire \epcs|readdata[14]~10_combout ;
wire \sdram|za_data[14]~q ;
wire \epcs|readdata[15]~11_combout ;
wire \sdram|za_data[15]~q ;
wire \epcs|readdata[10]~12_combout ;
wire \sdram|za_data[10]~q ;
wire \epcs|readdata[9]~13_combout ;
wire \sdram|za_data[9]~q ;
wire \epcs|readdata[8]~14_combout ;
wire \sdram|za_data[8]~q ;
wire \epcs|readdata[7]~15_combout ;
wire \sdram|za_data[7]~q ;
wire \epcs|readdata[6]~16_combout ;
wire \sdram|za_data[6]~q ;
wire \epcs|readdata[21]~17_combout ;
wire \epcs|readdata[30]~18_combout ;
wire \epcs|readdata[29]~19_combout ;
wire \epcs|readdata[28]~20_combout ;
wire \epcs|readdata[27]~21_combout ;
wire \epcs|readdata[26]~22_combout ;
wire \epcs|readdata[25]~23_combout ;
wire \epcs|readdata[24]~24_combout ;
wire \epcs|readdata[23]~25_combout ;
wire \epcs|readdata[22]~26_combout ;
wire \epcs|readdata[20]~27_combout ;
wire \epcs|readdata[19]~28_combout ;
wire \epcs|readdata[18]~29_combout ;
wire \epcs|readdata[17]~30_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~9_combout ;
wire \jtag|read_0~q ;
wire \jtag|av_readdata[0]~0_combout ;
wire \sys_pll|readdata[0]~1_combout ;
wire \epcs|the_niosII_epcs_sub|irq_reg~q ;
wire \jtag|av_readdata[9]~combout ;
wire \jtag|av_irq~combout ;
wire \rst_controller_001|r_early_rst~q ;
wire \mm_interconnect_0|cmd_mux_010|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_010|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_010|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_010|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_010|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~10_combout ;
wire \jtag|av_readdata[1]~1_combout ;
wire \sys_pll|readdata[1]~2_combout ;
wire \jtag|av_readdata[2]~2_combout ;
wire \jtag|av_readdata[3]~3_combout ;
wire \jtag|av_readdata[4]~4_combout ;
wire \jtag|av_readdata[5]~5_combout ;
wire \jtag|av_readdata[6]~6_combout ;
wire \jtag|av_readdata[7]~7_combout ;
wire \rs232_0|data_to_uart[4]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[2]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~13_combout ;
wire \epcs|readdata[31]~31_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~28_combout ;
wire \jtag|rvalid~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~29_combout ;
wire \jtag|woverflow~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~31_combout ;
wire \jtag|ac~q ;
wire \jtag|av_readdata[8]~8_combout ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[1]~q ;
wire \rs232_0|data_to_uart[5]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[3]~q ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~32_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_010|src_payload~17_combout ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[10]~q ;
wire \rs232_0|data_to_uart[6]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[4]~q ;
wire \rs232_0|data_to_uart[7]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[5]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[6]~q ;
wire \mm_interconnect_0|port_sw_avalon_parallel_port_slave_agent_rsp_fifo|write~3_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \port_gpio_0_export[0]~input_o ;
wire \port_gpio_0_export[1]~input_o ;
wire \port_gpio_0_export[2]~input_o ;
wire \port_gpio_0_export[3]~input_o ;
wire \port_gpio_0_export[4]~input_o ;
wire \port_gpio_0_export[5]~input_o ;
wire \port_gpio_0_export[6]~input_o ;
wire \port_gpio_0_export[7]~input_o ;
wire \port_gpio_0_export[8]~input_o ;
wire \port_gpio_0_export[9]~input_o ;
wire \port_gpio_0_export[10]~input_o ;
wire \port_gpio_0_export[11]~input_o ;
wire \port_gpio_0_export[12]~input_o ;
wire \port_gpio_0_export[13]~input_o ;
wire \port_gpio_0_export[14]~input_o ;
wire \port_gpio_0_export[15]~input_o ;
wire \port_gpio_0_export[16]~input_o ;
wire \port_gpio_0_export[17]~input_o ;
wire \port_gpio_0_export[18]~input_o ;
wire \port_gpio_0_export[19]~input_o ;
wire \port_gpio_0_export[20]~input_o ;
wire \port_gpio_0_export[21]~input_o ;
wire \port_gpio_0_export[22]~input_o ;
wire \port_gpio_0_export[23]~input_o ;
wire \port_gpio_0_export[24]~input_o ;
wire \port_gpio_0_export[25]~input_o ;
wire \port_gpio_0_export[26]~input_o ;
wire \port_gpio_0_export[27]~input_o ;
wire \port_gpio_0_export[28]~input_o ;
wire \port_gpio_0_export[29]~input_o ;
wire \port_gpio_0_export[30]~input_o ;
wire \port_gpio_0_export[31]~input_o ;
wire \sdram_dq[0]~input_o ;
wire \sdram_dq[1]~input_o ;
wire \sdram_dq[2]~input_o ;
wire \sdram_dq[3]~input_o ;
wire \sdram_dq[4]~input_o ;
wire \sdram_dq[5]~input_o ;
wire \sdram_dq[6]~input_o ;
wire \sdram_dq[7]~input_o ;
wire \sdram_dq[8]~input_o ;
wire \sdram_dq[9]~input_o ;
wire \sdram_dq[10]~input_o ;
wire \sdram_dq[11]~input_o ;
wire \sdram_dq[12]~input_o ;
wire \sdram_dq[13]~input_o ;
wire \sdram_dq[14]~input_o ;
wire \sdram_dq[15]~input_o ;
wire \clk_clk~input_o ;
wire \reset_reset_n~input_o ;
wire \port_sw_export[0]~input_o ;
wire \port_key_export[0]~input_o ;
wire \port_sw_export[1]~input_o ;
wire \port_key_export[1]~input_o ;
wire \port_sw_export[2]~input_o ;
wire \port_sw_export[3]~input_o ;
wire \adc_0_dout~input_o ;
wire \epcs_data0~input_o ;
wire \rs232_0_RXD~input_o ;
wire \rs232_1_RXD~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~8 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~16 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


niosII_niosII_epcs epcs(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.SCLK_reg(\epcs|the_niosII_epcs_sub|SCLK_reg~q ),
	.sce(\epcs|the_niosII_epcs_sub|SS_n~0_combout ),
	.shift_reg_7(\epcs|the_niosII_epcs_sub|shift_reg[7]~q ),
	.r_sync_rst(\rst_controller_001|r_sync_rst~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_010|saved_grant[0]~q ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_010|saved_grant[1]~q ),
	.out_data_buffer_38(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[38]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_010|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_010|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_010|src_data[40]~combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_010|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_010|src_payload~1_combout ),
	.mem_used_1(\mm_interconnect_0|epcs_epcs_control_port_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|epcs_epcs_control_port_translator|wait_latency_counter[1]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_010|src_valid~0_combout ),
	.src_valid1(\mm_interconnect_0|cmd_mux_010|src_valid~1_combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_010|src_data[46]~combout ),
	.out_data_buffer_65(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[65]~q ),
	.p1_wr_strobe(\epcs|the_niosII_epcs_sub|p1_wr_strobe~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_010|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_010|src_payload~3_combout ),
	.src_data_66(\mm_interconnect_0|cmd_mux_010|src_data[66]~combout ),
	.av_begintransfer(\mm_interconnect_0|epcs_epcs_control_port_translator|av_begintransfer~0_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_010|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_010|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_010|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_010|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_010|src_payload~8_combout ),
	.readdata_0(\epcs|readdata[0]~0_combout ),
	.readdata_1(\epcs|readdata[1]~1_combout ),
	.readdata_2(\epcs|readdata[2]~2_combout ),
	.readdata_3(\epcs|readdata[3]~3_combout ),
	.readdata_4(\epcs|readdata[4]~4_combout ),
	.readdata_11(\epcs|readdata[11]~5_combout ),
	.readdata_13(\epcs|readdata[13]~6_combout ),
	.readdata_16(\epcs|readdata[16]~7_combout ),
	.readdata_12(\epcs|readdata[12]~8_combout ),
	.readdata_5(\epcs|readdata[5]~9_combout ),
	.readdata_14(\epcs|readdata[14]~10_combout ),
	.readdata_15(\epcs|readdata[15]~11_combout ),
	.readdata_10(\epcs|readdata[10]~12_combout ),
	.readdata_9(\epcs|readdata[9]~13_combout ),
	.readdata_8(\epcs|readdata[8]~14_combout ),
	.readdata_7(\epcs|readdata[7]~15_combout ),
	.readdata_6(\epcs|readdata[6]~16_combout ),
	.readdata_21(\epcs|readdata[21]~17_combout ),
	.readdata_30(\epcs|readdata[30]~18_combout ),
	.readdata_29(\epcs|readdata[29]~19_combout ),
	.readdata_28(\epcs|readdata[28]~20_combout ),
	.readdata_27(\epcs|readdata[27]~21_combout ),
	.readdata_26(\epcs|readdata[26]~22_combout ),
	.readdata_25(\epcs|readdata[25]~23_combout ),
	.readdata_24(\epcs|readdata[24]~24_combout ),
	.readdata_23(\epcs|readdata[23]~25_combout ),
	.readdata_22(\epcs|readdata[22]~26_combout ),
	.readdata_20(\epcs|readdata[20]~27_combout ),
	.readdata_19(\epcs|readdata[19]~28_combout ),
	.readdata_18(\epcs|readdata[18]~29_combout ),
	.readdata_17(\epcs|readdata[17]~30_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_010|src_payload~9_combout ),
	.irq_reg(\epcs|the_niosII_epcs_sub|irq_reg~q ),
	.r_early_rst(\rst_controller_001|r_early_rst~q ),
	.src_data_41(\mm_interconnect_0|cmd_mux_010|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_010|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_010|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_010|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_010|src_data[45]~combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_010|src_payload~10_combout ),
	.readdata_31(\epcs|readdata[31]~31_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_010|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_010|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_010|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_010|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_010|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_010|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_010|src_payload~17_combout ),
	.epcs_data0(\epcs_data0~input_o ));

niosII_niosII_jtag jtag(
	.tdo(\jtag|niosII_jtag_alt_jtag_atlantic|tdo~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.rst1(\jtag|niosII_jtag_alt_jtag_atlantic|rst1~q ),
	.b_full(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.out_data_toggle_flopped(\mm_interconnect_0|crosser|clock_xer|out_data_toggle_flopped~q ),
	.b_non_empty(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_5(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.dreg_0(\mm_interconnect_0|crosser|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.av_waitrequest1(\jtag|av_waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|jtag_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.out_data_buffer_66(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[66]~q ),
	.out_data_buffer_38(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_7(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[7]~q ),
	.out_data_buffer_65(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[65]~q ),
	.out_data_buffer_0(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[0]~q ),
	.b_full1(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_21(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_11(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_51(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_41(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_31(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_01(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.out_data_buffer_1(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[1]~q ),
	.read_01(\jtag|read_0~q ),
	.av_readdata_0(\jtag|av_readdata[0]~0_combout ),
	.av_readdata_9(\jtag|av_readdata[9]~combout ),
	.av_irq1(\jtag|av_irq~combout ),
	.av_readdata_1(\jtag|av_readdata[1]~1_combout ),
	.av_readdata_2(\jtag|av_readdata[2]~2_combout ),
	.av_readdata_3(\jtag|av_readdata[3]~3_combout ),
	.av_readdata_4(\jtag|av_readdata[4]~4_combout ),
	.av_readdata_5(\jtag|av_readdata[5]~5_combout ),
	.av_readdata_6(\jtag|av_readdata[6]~6_combout ),
	.av_readdata_7(\jtag|av_readdata[7]~7_combout ),
	.out_data_buffer_2(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[2]~q ),
	.rvalid1(\jtag|rvalid~q ),
	.woverflow1(\jtag|woverflow~q ),
	.ac1(\jtag|ac~q ),
	.av_readdata_8(\jtag|av_readdata[8]~8_combout ),
	.out_data_buffer_3(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_10(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_4(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_5(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_6(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[6]~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

niosII_niosII_rs232_0 rs232_0(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.readdata_0(\rs232_0|readdata[0]~q ),
	.irq1(\rs232_0|irq~q ),
	.readdata_1(\rs232_0|readdata[1]~q ),
	.readdata_23(\rs232_0|readdata[23]~q ),
	.readdata_22(\rs232_0|readdata[22]~q ),
	.readdata_21(\rs232_0|readdata[21]~q ),
	.readdata_20(\rs232_0|readdata[20]~q ),
	.readdata_19(\rs232_0|readdata[19]~q ),
	.readdata_18(\rs232_0|readdata[18]~q ),
	.readdata_17(\rs232_0|readdata[17]~q ),
	.readdata_16(\rs232_0|readdata[16]~q ),
	.serial_data_out(\rs232_0|RS232_Out_Serializer|serial_data_out~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_read(\cpu|cpu|d_read~q ),
	.read_accepted(\mm_interconnect_0|cpu_data_master_translator|read_accepted~q ),
	.hold_waitrequest(\mm_interconnect_0|cpu_data_master_agent|hold_waitrequest~q ),
	.cp_valid(\mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ),
	.data(\port_led|data~0_combout ),
	.d_byteenable_0(\cpu|cpu|d_byteenable[0]~q ),
	.Equal9(\mm_interconnect_0|router|Equal9~0_combout ),
	.data1(\port_led|data~3_combout ),
	.data2(\port_led|data~4_combout ),
	.data3(\port_led|data~5_combout ),
	.data4(\port_led|data~6_combout ),
	.data5(\port_led|data~7_combout ),
	.data6(\port_led|data~8_combout ),
	.data7(\port_led|data~9_combout ),
	.Equal12(\mm_interconnect_0|router|Equal12~1_combout ),
	.mem_used_1(\mm_interconnect_0|rs232_0_avalon_rs232_slave_agent_rsp_fifo|mem_used[1]~q ),
	.Equal121(\mm_interconnect_0|router|Equal12~2_combout ),
	.data_to_uart_0(\rs232_0|data_to_uart[0]~q ),
	.data8(\port_led|data~10_combout ),
	.read_latency_shift_reg(\mm_interconnect_0|rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg~1_combout ),
	.readdata_2(\rs232_0|readdata[2]~q ),
	.readdata_3(\rs232_0|readdata[3]~q ),
	.readdata_4(\rs232_0|readdata[4]~q ),
	.readdata_5(\rs232_0|readdata[5]~q ),
	.readdata_6(\rs232_0|readdata[6]~q ),
	.readdata_7(\rs232_0|readdata[7]~q ),
	.data_to_uart_1(\rs232_0|data_to_uart[1]~q ),
	.readdata_15(\rs232_0|readdata[15]~q ),
	.readdata_9(\rs232_0|readdata[9]~q ),
	.readdata_8(\rs232_0|readdata[8]~q ),
	.data_to_uart_2(\rs232_0|data_to_uart[2]~q ),
	.comb(\rs232_0|RS232_In_Deserializer|comb~1_combout ),
	.data_to_uart_3(\rs232_0|data_to_uart[3]~q ),
	.data_to_uart_4(\rs232_0|data_to_uart[4]~q ),
	.data_to_uart_5(\rs232_0|data_to_uart[5]~q ),
	.data_to_uart_6(\rs232_0|data_to_uart[6]~q ),
	.data_to_uart_7(\rs232_0|data_to_uart[7]~q ),
	.GND_port(\~GND~combout ),
	.rs232_0_RXD(\rs232_0_RXD~input_o ));

niosII_niosII_port_sw port_sw(
	.clk(\sys_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.cp_valid(\mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ),
	.write(\mm_interconnect_0|port_sw_avalon_parallel_port_slave_agent_rsp_fifo|write~2_combout ),
	.readdata_0(\port_sw|readdata[0]~q ),
	.readdata_1(\port_sw|readdata[1]~q ),
	.readdata_2(\port_sw|readdata[2]~q ),
	.readdata_3(\port_sw|readdata[3]~q ),
	.DIP({\port_sw_export[3]~input_o ,\port_sw_export[2]~input_o ,\port_sw_export[1]~input_o ,\port_sw_export[0]~input_o }));

niosII_niosII_port_led port_led(
	.clk(\sys_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.data_out_0(\port_led|data_out[0]~q ),
	.data_out_1(\port_led|data_out[1]~q ),
	.data_out_2(\port_led|data_out[2]~q ),
	.data_out_3(\port_led|data_out[3]~q ),
	.data_out_4(\port_led|data_out[4]~q ),
	.data_out_5(\port_led|data_out[5]~q ),
	.data_out_6(\port_led|data_out[6]~q ),
	.data_out_7(\port_led|data_out[7]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.hold_waitrequest(\mm_interconnect_0|cpu_data_master_agent|hold_waitrequest~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|cpu_data_master_translator|write_accepted~q ),
	.cp_valid(\mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ),
	.d_writedata_0(\cpu|cpu|d_writedata[0]~q ),
	.data(\port_led|data~0_combout ),
	.d_byteenable_0(\cpu|cpu|d_byteenable[0]~q ),
	.Equal6(\timer_0|Equal6~0_combout ),
	.read_latency_shift_reg(\mm_interconnect_0|port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg~0_combout ),
	.d_writedata_1(\cpu|cpu|d_writedata[1]~q ),
	.data1(\port_led|data~3_combout ),
	.d_writedata_2(\cpu|cpu|d_writedata[2]~q ),
	.data2(\port_led|data~4_combout ),
	.d_writedata_3(\cpu|cpu|d_writedata[3]~q ),
	.data3(\port_led|data~5_combout ),
	.d_writedata_4(\cpu|cpu|d_writedata[4]~q ),
	.data4(\port_led|data~6_combout ),
	.d_writedata_5(\cpu|cpu|d_writedata[5]~q ),
	.data5(\port_led|data~7_combout ),
	.d_writedata_6(\cpu|cpu|d_writedata[6]~q ),
	.data6(\port_led|data~8_combout ),
	.d_writedata_7(\cpu|cpu|d_writedata[7]~q ),
	.data7(\port_led|data~9_combout ),
	.data8(\port_led|data~10_combout ),
	.readdata_0(\port_led|readdata[0]~q ),
	.readdata_1(\port_led|readdata[1]~q ),
	.readdata_2(\port_led|readdata[2]~q ),
	.readdata_3(\port_led|readdata[3]~q ),
	.readdata_4(\port_led|readdata[4]~q ),
	.readdata_5(\port_led|readdata[5]~q ),
	.readdata_6(\port_led|readdata[6]~q ),
	.readdata_7(\port_led|readdata[7]~q ));

niosII_niosII_port_key port_key(
	.clk(\sys_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.cp_valid(\mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ),
	.write(\mm_interconnect_0|port_key_avalon_parallel_port_slave_agent_rsp_fifo|write~0_combout ),
	.readdata_0(\port_key|readdata[0]~q ),
	.readdata_1(\port_key|readdata[1]~q ),
	.port_key_export_0(\port_key_export[0]~input_o ),
	.port_key_export_1(\port_key_export[1]~input_o ));

niosII_niosII_port_gpio_0 port_gpio_0(
	.clk(\sys_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.d_writedata_24(\cpu|cpu|d_writedata[24]~q ),
	.d_writedata_25(\cpu|cpu|d_writedata[25]~q ),
	.d_writedata_26(\cpu|cpu|d_writedata[26]~q ),
	.d_writedata_27(\cpu|cpu|d_writedata[27]~q ),
	.d_writedata_28(\cpu|cpu|d_writedata[28]~q ),
	.d_writedata_29(\cpu|cpu|d_writedata[29]~q ),
	.d_writedata_30(\cpu|cpu|d_writedata[30]~q ),
	.d_writedata_31(\cpu|cpu|d_writedata[31]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.cp_valid(\mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ),
	.m0_write(\mm_interconnect_0|timer_0_s1_agent|m0_write~0_combout ),
	.data(\port_led|data~0_combout ),
	.d_byteenable_0(\cpu|cpu|d_byteenable[0]~q ),
	.data1(\port_led|data~3_combout ),
	.data2(\port_led|data~4_combout ),
	.data3(\port_led|data~5_combout ),
	.data4(\port_led|data~6_combout ),
	.data5(\port_led|data~7_combout ),
	.data6(\port_led|data~8_combout ),
	.data7(\port_led|data~9_combout ),
	.d_byteenable_1(\cpu|cpu|d_byteenable[1]~q ),
	.data_out_0(\port_gpio_0|data_out[0]~q ),
	.direction_0(\port_gpio_0|direction[0]~q ),
	.data_out_1(\port_gpio_0|data_out[1]~q ),
	.direction_1(\port_gpio_0|direction[1]~q ),
	.data_out_2(\port_gpio_0|data_out[2]~q ),
	.direction_2(\port_gpio_0|direction[2]~q ),
	.data_out_3(\port_gpio_0|data_out[3]~q ),
	.direction_3(\port_gpio_0|direction[3]~q ),
	.data_out_4(\port_gpio_0|data_out[4]~q ),
	.direction_4(\port_gpio_0|direction[4]~q ),
	.data_out_5(\port_gpio_0|data_out[5]~q ),
	.direction_5(\port_gpio_0|direction[5]~q ),
	.data_out_6(\port_gpio_0|data_out[6]~q ),
	.direction_6(\port_gpio_0|direction[6]~q ),
	.data_out_7(\port_gpio_0|data_out[7]~q ),
	.direction_7(\port_gpio_0|direction[7]~q ),
	.data_out_8(\port_gpio_0|data_out[8]~q ),
	.direction_8(\port_gpio_0|direction[8]~q ),
	.data_out_9(\port_gpio_0|data_out[9]~q ),
	.direction_9(\port_gpio_0|direction[9]~q ),
	.data_out_10(\port_gpio_0|data_out[10]~q ),
	.direction_10(\port_gpio_0|direction[10]~q ),
	.data_out_11(\port_gpio_0|data_out[11]~q ),
	.direction_11(\port_gpio_0|direction[11]~q ),
	.data_out_12(\port_gpio_0|data_out[12]~q ),
	.direction_12(\port_gpio_0|direction[12]~q ),
	.data_out_13(\port_gpio_0|data_out[13]~q ),
	.direction_13(\port_gpio_0|direction[13]~q ),
	.data_out_14(\port_gpio_0|data_out[14]~q ),
	.direction_14(\port_gpio_0|direction[14]~q ),
	.data_out_15(\port_gpio_0|data_out[15]~q ),
	.direction_15(\port_gpio_0|direction[15]~q ),
	.data_out_16(\port_gpio_0|data_out[16]~q ),
	.direction_16(\port_gpio_0|direction[16]~q ),
	.data_out_17(\port_gpio_0|data_out[17]~q ),
	.direction_17(\port_gpio_0|direction[17]~q ),
	.data_out_18(\port_gpio_0|data_out[18]~q ),
	.direction_18(\port_gpio_0|direction[18]~q ),
	.data_out_19(\port_gpio_0|data_out[19]~q ),
	.direction_19(\port_gpio_0|direction[19]~q ),
	.data_out_20(\port_gpio_0|data_out[20]~q ),
	.direction_20(\port_gpio_0|direction[20]~q ),
	.data_out_21(\port_gpio_0|data_out[21]~q ),
	.direction_21(\port_gpio_0|direction[21]~q ),
	.data_out_22(\port_gpio_0|data_out[22]~q ),
	.direction_22(\port_gpio_0|direction[22]~q ),
	.data_out_23(\port_gpio_0|data_out[23]~q ),
	.direction_23(\port_gpio_0|direction[23]~q ),
	.data_out_24(\port_gpio_0|data_out[24]~q ),
	.direction_24(\port_gpio_0|direction[24]~q ),
	.data_out_25(\port_gpio_0|data_out[25]~q ),
	.direction_25(\port_gpio_0|direction[25]~q ),
	.data_out_26(\port_gpio_0|data_out[26]~q ),
	.direction_26(\port_gpio_0|direction[26]~q ),
	.data_out_27(\port_gpio_0|data_out[27]~q ),
	.direction_27(\port_gpio_0|direction[27]~q ),
	.data_out_28(\port_gpio_0|data_out[28]~q ),
	.direction_28(\port_gpio_0|direction[28]~q ),
	.data_out_29(\port_gpio_0|data_out[29]~q ),
	.direction_29(\port_gpio_0|direction[29]~q ),
	.data_out_30(\port_gpio_0|data_out[30]~q ),
	.direction_30(\port_gpio_0|direction[30]~q ),
	.data_out_31(\port_gpio_0|data_out[31]~q ),
	.direction_31(\port_gpio_0|direction[31]~q ),
	.d_writedata_10(\cpu|cpu|d_writedata[10]~q ),
	.d_byteenable_2(\cpu|cpu|d_byteenable[2]~q ),
	.d_byteenable_3(\cpu|cpu|d_byteenable[3]~q ),
	.read_latency_shift_reg(\mm_interconnect_0|port_gpio_0_avalon_parallel_port_slave_translator|read_latency_shift_reg~0_combout ),
	.d_writedata_8(\cpu|cpu|d_writedata[8]~q ),
	.d_writedata_9(\cpu|cpu|d_writedata[9]~q ),
	.d_writedata_11(\cpu|cpu|d_writedata[11]~q ),
	.d_writedata_12(\cpu|cpu|d_writedata[12]~q ),
	.d_writedata_13(\cpu|cpu|d_writedata[13]~q ),
	.d_writedata_14(\cpu|cpu|d_writedata[14]~q ),
	.d_writedata_15(\cpu|cpu|d_writedata[15]~q ),
	.d_writedata_16(\cpu|cpu|d_writedata[16]~q ),
	.d_writedata_17(\cpu|cpu|d_writedata[17]~q ),
	.d_writedata_18(\cpu|cpu|d_writedata[18]~q ),
	.d_writedata_19(\cpu|cpu|d_writedata[19]~q ),
	.d_writedata_20(\cpu|cpu|d_writedata[20]~q ),
	.d_writedata_21(\cpu|cpu|d_writedata[21]~q ),
	.d_writedata_22(\cpu|cpu|d_writedata[22]~q ),
	.d_writedata_23(\cpu|cpu|d_writedata[23]~q ),
	.readdata_0(\port_gpio_0|readdata[0]~q ),
	.readdata_1(\port_gpio_0|readdata[1]~q ),
	.readdata_2(\port_gpio_0|readdata[2]~q ),
	.readdata_3(\port_gpio_0|readdata[3]~q ),
	.readdata_4(\port_gpio_0|readdata[4]~q ),
	.readdata_5(\port_gpio_0|readdata[5]~q ),
	.readdata_6(\port_gpio_0|readdata[6]~q ),
	.readdata_7(\port_gpio_0|readdata[7]~q ),
	.readdata_26(\port_gpio_0|readdata[26]~q ),
	.readdata_25(\port_gpio_0|readdata[25]~q ),
	.readdata_24(\port_gpio_0|readdata[24]~q ),
	.readdata_23(\port_gpio_0|readdata[23]~q ),
	.readdata_22(\port_gpio_0|readdata[22]~q ),
	.readdata_21(\port_gpio_0|readdata[21]~q ),
	.readdata_20(\port_gpio_0|readdata[20]~q ),
	.readdata_19(\port_gpio_0|readdata[19]~q ),
	.readdata_18(\port_gpio_0|readdata[18]~q ),
	.readdata_17(\port_gpio_0|readdata[17]~q ),
	.readdata_16(\port_gpio_0|readdata[16]~q ),
	.readdata_15(\port_gpio_0|readdata[15]~q ),
	.readdata_14(\port_gpio_0|readdata[14]~q ),
	.readdata_13(\port_gpio_0|readdata[13]~q ),
	.readdata_12(\port_gpio_0|readdata[12]~q ),
	.readdata_11(\port_gpio_0|readdata[11]~q ),
	.readdata_10(\port_gpio_0|readdata[10]~q ),
	.readdata_9(\port_gpio_0|readdata[9]~q ),
	.readdata_8(\port_gpio_0|readdata[8]~q ),
	.readdata_27(\port_gpio_0|readdata[27]~q ),
	.readdata_28(\port_gpio_0|readdata[28]~q ),
	.readdata_29(\port_gpio_0|readdata[29]~q ),
	.readdata_30(\port_gpio_0|readdata[30]~q ),
	.readdata_31(\port_gpio_0|readdata[31]~q ),
	.port_gpio_0_export_0(\port_gpio_0_export[0]~input_o ),
	.port_gpio_0_export_1(\port_gpio_0_export[1]~input_o ),
	.port_gpio_0_export_2(\port_gpio_0_export[2]~input_o ),
	.port_gpio_0_export_3(\port_gpio_0_export[3]~input_o ),
	.port_gpio_0_export_4(\port_gpio_0_export[4]~input_o ),
	.port_gpio_0_export_5(\port_gpio_0_export[5]~input_o ),
	.port_gpio_0_export_6(\port_gpio_0_export[6]~input_o ),
	.port_gpio_0_export_7(\port_gpio_0_export[7]~input_o ),
	.port_gpio_0_export_8(\port_gpio_0_export[8]~input_o ),
	.port_gpio_0_export_9(\port_gpio_0_export[9]~input_o ),
	.port_gpio_0_export_10(\port_gpio_0_export[10]~input_o ),
	.port_gpio_0_export_11(\port_gpio_0_export[11]~input_o ),
	.port_gpio_0_export_12(\port_gpio_0_export[12]~input_o ),
	.port_gpio_0_export_13(\port_gpio_0_export[13]~input_o ),
	.port_gpio_0_export_14(\port_gpio_0_export[14]~input_o ),
	.port_gpio_0_export_15(\port_gpio_0_export[15]~input_o ),
	.port_gpio_0_export_16(\port_gpio_0_export[16]~input_o ),
	.port_gpio_0_export_17(\port_gpio_0_export[17]~input_o ),
	.port_gpio_0_export_18(\port_gpio_0_export[18]~input_o ),
	.port_gpio_0_export_19(\port_gpio_0_export[19]~input_o ),
	.port_gpio_0_export_20(\port_gpio_0_export[20]~input_o ),
	.port_gpio_0_export_21(\port_gpio_0_export[21]~input_o ),
	.port_gpio_0_export_22(\port_gpio_0_export[22]~input_o ),
	.port_gpio_0_export_23(\port_gpio_0_export[23]~input_o ),
	.port_gpio_0_export_24(\port_gpio_0_export[24]~input_o ),
	.port_gpio_0_export_25(\port_gpio_0_export[25]~input_o ),
	.port_gpio_0_export_26(\port_gpio_0_export[26]~input_o ),
	.port_gpio_0_export_27(\port_gpio_0_export[27]~input_o ),
	.port_gpio_0_export_28(\port_gpio_0_export[28]~input_o ),
	.port_gpio_0_export_29(\port_gpio_0_export[29]~input_o ),
	.port_gpio_0_export_30(\port_gpio_0_export[30]~input_o ),
	.port_gpio_0_export_31(\port_gpio_0_export[31]~input_o ));

niosII_niosII_rs232_0_1 rs232_1(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.readdata_0(\rs232_1|readdata[0]~q ),
	.irq1(\rs232_1|irq~q ),
	.readdata_1(\rs232_1|readdata[1]~q ),
	.readdata_23(\rs232_1|readdata[23]~q ),
	.readdata_22(\rs232_1|readdata[22]~q ),
	.readdata_21(\rs232_1|readdata[21]~q ),
	.readdata_20(\rs232_1|readdata[20]~q ),
	.readdata_19(\rs232_1|readdata[19]~q ),
	.readdata_18(\rs232_1|readdata[18]~q ),
	.readdata_17(\rs232_1|readdata[17]~q ),
	.readdata_16(\rs232_1|readdata[16]~q ),
	.serial_data_out(\rs232_1|RS232_Out_Serializer|serial_data_out~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.cp_valid(\mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ),
	.data(\port_led|data~0_combout ),
	.data1(\port_led|data~3_combout ),
	.read_latency_shift_reg(\mm_interconnect_0|rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg~2_combout ),
	.data_to_uart_0(\rs232_0|data_to_uart[0]~q ),
	.data2(\port_led|data~10_combout ),
	.readdata_2(\rs232_1|readdata[2]~q ),
	.readdata_3(\rs232_1|readdata[3]~q ),
	.readdata_4(\rs232_1|readdata[4]~q ),
	.readdata_5(\rs232_1|readdata[5]~q ),
	.readdata_6(\rs232_1|readdata[6]~q ),
	.readdata_7(\rs232_1|readdata[7]~q ),
	.data_to_uart_1(\rs232_0|data_to_uart[1]~q ),
	.readdata_15(\rs232_1|readdata[15]~q ),
	.readdata_9(\rs232_1|readdata[9]~q ),
	.readdata_8(\rs232_1|readdata[8]~q ),
	.data_to_uart_2(\rs232_0|data_to_uart[2]~q ),
	.comb(\rs232_0|RS232_In_Deserializer|comb~1_combout ),
	.data_to_uart_3(\rs232_0|data_to_uart[3]~q ),
	.data_to_uart_4(\rs232_0|data_to_uart[4]~q ),
	.data_to_uart_5(\rs232_0|data_to_uart[5]~q ),
	.data_to_uart_6(\rs232_0|data_to_uart[6]~q ),
	.data_to_uart_7(\rs232_0|data_to_uart[7]~q ),
	.GND_port(\~GND~combout ),
	.rs232_1_RXD(\rs232_1_RXD~input_o ));

niosII_niosII_sdram sdram(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.m_addr_0(\sdram|m_addr[0]~q ),
	.m_addr_1(\sdram|m_addr[1]~q ),
	.m_addr_2(\sdram|m_addr[2]~q ),
	.m_addr_3(\sdram|m_addr[3]~q ),
	.m_addr_4(\sdram|m_addr[4]~q ),
	.m_addr_5(\sdram|m_addr[5]~q ),
	.m_addr_6(\sdram|m_addr[6]~q ),
	.m_addr_7(\sdram|m_addr[7]~q ),
	.m_addr_8(\sdram|m_addr[8]~q ),
	.byteen_reg_0(\mm_interconnect_0|sdram_s1_cmd_width_adapter|byteen_reg[0]~q ),
	.byteen_reg_1(\mm_interconnect_0|sdram_s1_cmd_width_adapter|byteen_reg[1]~q ),
	.oe1(\sdram|oe~q ),
	.m_addr_9(\sdram|m_addr[9]~q ),
	.m_addr_10(\sdram|m_addr[10]~q ),
	.m_addr_11(\sdram|m_addr[11]~q ),
	.m_addr_12(\sdram|m_addr[12]~q ),
	.m_bank_0(\sdram|m_bank[0]~q ),
	.m_bank_1(\sdram|m_bank[1]~q ),
	.m_cmd_1(\sdram|m_cmd[1]~q ),
	.m_cmd_3(\sdram|m_cmd[3]~q ),
	.m_dqm_0(\sdram|m_dqm[0]~q ),
	.m_dqm_1(\sdram|m_dqm[1]~q ),
	.m_cmd_2(\sdram|m_cmd[2]~q ),
	.m_cmd_0(\sdram|m_cmd[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.entries_1(\sdram|the_niosII_sdram_input_efifo_module|entries[1]~q ),
	.entries_0(\sdram|the_niosII_sdram_input_efifo_module|entries[0]~q ),
	.d_byteenable_0(\cpu|cpu|d_byteenable[0]~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_012|saved_grant[0]~q ),
	.d_byteenable_1(\cpu|cpu|d_byteenable[1]~q ),
	.use_reg(\mm_interconnect_0|sdram_s1_cmd_width_adapter|use_reg~q ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_012|saved_grant[1]~q ),
	.WideOr0(\mm_interconnect_0|sdram_s1_agent|WideOr0~2_combout ),
	.Equal0(\sdram|the_niosII_sdram_input_efifo_module|Equal0~0_combout ),
	.Equal1(\mm_interconnect_0|router|Equal1~0_combout ),
	.WideOr1(\mm_interconnect_0|cmd_mux_012|WideOr1~combout ),
	.m0_write(\mm_interconnect_0|sdram_s1_agent|m0_write~2_combout ),
	.mem_used_7(\mm_interconnect_0|sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.src_data_66(\mm_interconnect_0|cmd_mux_012|src_data[66]~combout ),
	.out_data_28(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[28]~0_combout ),
	.src_valid(\mm_interconnect_0|cmd_mux_012|src_valid~0_combout ),
	.src12_valid(\mm_interconnect_0|cmd_demux|src12_valid~0_combout ),
	.m0_write1(\mm_interconnect_0|sdram_s1_agent|m0_write~combout ),
	.out_data_42(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[42]~1_combout ),
	.out_data_29(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[29]~2_combout ),
	.out_data_31(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[31]~3_combout ),
	.out_data_30(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[30]~4_combout ),
	.out_data_33(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[33]~5_combout ),
	.out_data_32(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[32]~6_combout ),
	.out_data_35(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[35]~7_combout ),
	.out_data_34(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[34]~8_combout ),
	.out_data_37(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[37]~9_combout ),
	.out_data_36(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[36]~10_combout ),
	.out_data_39(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[39]~11_combout ),
	.out_data_38(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[38]~12_combout ),
	.out_data_41(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[41]~13_combout ),
	.out_data_40(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[40]~14_combout ),
	.out_data_19(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[19]~15_combout ),
	.out_data_20(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[20]~16_combout ),
	.out_data_21(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[21]~17_combout ),
	.out_data_22(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[22]~18_combout ),
	.out_data_23(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[23]~19_combout ),
	.out_data_24(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[24]~20_combout ),
	.out_data_25(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[25]~21_combout ),
	.out_data_26(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[26]~22_combout ),
	.out_data_27(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[27]~23_combout ),
	.m_data_0(\sdram|m_data[0]~q ),
	.m_data_1(\sdram|m_data[1]~q ),
	.m_data_2(\sdram|m_data[2]~q ),
	.m_data_3(\sdram|m_data[3]~q ),
	.m_data_4(\sdram|m_data[4]~q ),
	.m_data_5(\sdram|m_data[5]~q ),
	.m_data_6(\sdram|m_data[6]~q ),
	.m_data_7(\sdram|m_data[7]~q ),
	.m_data_8(\sdram|m_data[8]~q ),
	.m_data_9(\sdram|m_data[9]~q ),
	.m_data_10(\sdram|m_data[10]~q ),
	.m_data_11(\sdram|m_data[11]~q ),
	.m_data_12(\sdram|m_data[12]~q ),
	.m_data_13(\sdram|m_data[13]~q ),
	.m_data_14(\sdram|m_data[14]~q ),
	.m_data_15(\sdram|m_data[15]~q ),
	.out_data_0(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[0]~24_combout ),
	.out_data_1(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[1]~25_combout ),
	.out_data_2(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[2]~26_combout ),
	.out_data_3(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[3]~27_combout ),
	.out_data_4(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[4]~28_combout ),
	.out_data_5(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[5]~29_combout ),
	.out_data_6(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[6]~30_combout ),
	.out_data_7(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[7]~31_combout ),
	.out_data_8(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[8]~32_combout ),
	.out_data_9(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[9]~33_combout ),
	.out_data_10(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[10]~34_combout ),
	.out_data_11(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[11]~35_combout ),
	.out_data_12(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[12]~36_combout ),
	.out_data_13(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[13]~37_combout ),
	.out_data_14(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[14]~38_combout ),
	.out_data_15(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[15]~39_combout ),
	.za_valid1(\sdram|za_valid~q ),
	.za_data_0(\sdram|za_data[0]~q ),
	.za_data_1(\sdram|za_data[1]~q ),
	.za_data_2(\sdram|za_data[2]~q ),
	.za_data_3(\sdram|za_data[3]~q ),
	.za_data_4(\sdram|za_data[4]~q ),
	.za_data_11(\sdram|za_data[11]~q ),
	.za_data_13(\sdram|za_data[13]~q ),
	.za_data_12(\sdram|za_data[12]~q ),
	.za_data_5(\sdram|za_data[5]~q ),
	.za_data_14(\sdram|za_data[14]~q ),
	.za_data_15(\sdram|za_data[15]~q ),
	.za_data_10(\sdram|za_data[10]~q ),
	.za_data_9(\sdram|za_data[9]~q ),
	.za_data_8(\sdram|za_data[8]~q ),
	.za_data_7(\sdram|za_data[7]~q ),
	.za_data_6(\sdram|za_data[6]~q ),
	.sdram_dq_0(\sdram_dq[0]~input_o ),
	.sdram_dq_1(\sdram_dq[1]~input_o ),
	.sdram_dq_2(\sdram_dq[2]~input_o ),
	.sdram_dq_3(\sdram_dq[3]~input_o ),
	.sdram_dq_4(\sdram_dq[4]~input_o ),
	.sdram_dq_5(\sdram_dq[5]~input_o ),
	.sdram_dq_6(\sdram_dq[6]~input_o ),
	.sdram_dq_7(\sdram_dq[7]~input_o ),
	.sdram_dq_8(\sdram_dq[8]~input_o ),
	.sdram_dq_9(\sdram_dq[9]~input_o ),
	.sdram_dq_10(\sdram_dq[10]~input_o ),
	.sdram_dq_11(\sdram_dq[11]~input_o ),
	.sdram_dq_12(\sdram_dq[12]~input_o ),
	.sdram_dq_13(\sdram_dq[13]~input_o ),
	.sdram_dq_14(\sdram_dq[14]~input_o ),
	.sdram_dq_15(\sdram_dq[15]~input_o ));

niosII_niosII_mm_interconnect_0 mm_interconnect_0(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_6(\cpu|cpu|W_alu_result[6]~q ),
	.W_alu_result_26(\cpu|cpu|W_alu_result[26]~q ),
	.W_alu_result_25(\cpu|cpu|W_alu_result[25]~q ),
	.W_alu_result_24(\cpu|cpu|W_alu_result[24]~q ),
	.W_alu_result_23(\cpu|cpu|W_alu_result[23]~q ),
	.W_alu_result_22(\cpu|cpu|W_alu_result[22]~q ),
	.W_alu_result_21(\cpu|cpu|W_alu_result[21]~q ),
	.W_alu_result_20(\cpu|cpu|W_alu_result[20]~q ),
	.W_alu_result_19(\cpu|cpu|W_alu_result[19]~q ),
	.W_alu_result_18(\cpu|cpu|W_alu_result[18]~q ),
	.W_alu_result_17(\cpu|cpu|W_alu_result[17]~q ),
	.W_alu_result_16(\cpu|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\cpu|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\cpu|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\cpu|cpu|W_alu_result[13]~q ),
	.W_alu_result_12(\cpu|cpu|W_alu_result[12]~q ),
	.W_alu_result_11(\cpu|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\cpu|cpu|W_alu_result[10]~q ),
	.W_alu_result_5(\cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_7(\cpu|cpu|W_alu_result[7]~q ),
	.W_alu_result_9(\cpu|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\cpu|cpu|W_alu_result[8]~q ),
	.W_alu_result_4(\cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.byteen_reg_0(\mm_interconnect_0|sdram_s1_cmd_width_adapter|byteen_reg[0]~q ),
	.byteen_reg_1(\mm_interconnect_0|sdram_s1_cmd_width_adapter|byteen_reg[1]~q ),
	.d_writedata_24(\cpu|cpu|d_writedata[24]~q ),
	.d_writedata_25(\cpu|cpu|d_writedata[25]~q ),
	.d_writedata_26(\cpu|cpu|d_writedata[26]~q ),
	.d_writedata_27(\cpu|cpu|d_writedata[27]~q ),
	.d_writedata_28(\cpu|cpu|d_writedata[28]~q ),
	.d_writedata_29(\cpu|cpu|d_writedata[29]~q ),
	.d_writedata_30(\cpu|cpu|d_writedata[30]~q ),
	.d_writedata_31(\cpu|cpu|d_writedata[31]~q ),
	.readdata_0(\rs232_0|readdata[0]~q ),
	.readdata_01(\rs232_1|readdata[0]~q ),
	.readdata_4(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[4]~q ),
	.readdata_1(\rs232_0|readdata[1]~q ),
	.readdata_11(\rs232_1|readdata[1]~q ),
	.readdata_23(\rs232_0|readdata[23]~q ),
	.readdata_231(\rs232_1|readdata[23]~q ),
	.readdata_22(\rs232_1|readdata[22]~q ),
	.readdata_221(\rs232_0|readdata[22]~q ),
	.readdata_21(\rs232_1|readdata[21]~q ),
	.readdata_211(\rs232_0|readdata[21]~q ),
	.readdata_20(\rs232_1|readdata[20]~q ),
	.readdata_201(\rs232_0|readdata[20]~q ),
	.readdata_19(\rs232_1|readdata[19]~q ),
	.readdata_191(\rs232_0|readdata[19]~q ),
	.readdata_18(\rs232_1|readdata[18]~q ),
	.readdata_181(\rs232_0|readdata[18]~q ),
	.readdata_17(\rs232_1|readdata[17]~q ),
	.readdata_171(\rs232_0|readdata[17]~q ),
	.readdata_16(\rs232_1|readdata[16]~q ),
	.readdata_161(\rs232_0|readdata[16]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.r_sync_rst1(\rst_controller_001|r_sync_rst~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_010|saved_grant[0]~q ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_010|saved_grant[1]~q ),
	.out_data_buffer_38(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[38]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_010|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_010|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_010|src_data[40]~combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_010|src_payload~0_combout ),
	.entries_1(\sdram|the_niosII_sdram_input_efifo_module|entries[1]~q ),
	.entries_0(\sdram|the_niosII_sdram_input_efifo_module|entries[0]~q ),
	.mem_used_1(\mm_interconnect_0|adc_0_adc_slave_agent_rsp_fifo|mem_used[1]~q ),
	.d_read(\cpu|cpu|d_read~q ),
	.read_accepted(\mm_interconnect_0|cpu_data_master_translator|read_accepted~q ),
	.hold_waitrequest(\mm_interconnect_0|cpu_data_master_agent|hold_waitrequest~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|cpu_data_master_translator|write_accepted~q ),
	.cp_valid(\mm_interconnect_0|cpu_data_master_agent|cp_valid~0_combout ),
	.Equal3(\mm_interconnect_0|router|Equal3~6_combout ),
	.m0_read(\mm_interconnect_0|adc_0_adc_slave_agent|m0_read~combout ),
	.m0_write(\mm_interconnect_0|timer_0_s1_agent|m0_write~0_combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_010|src_payload~1_combout ),
	.mem_used_11(\mm_interconnect_0|epcs_epcs_control_port_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|epcs_epcs_control_port_translator|wait_latency_counter[1]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_010|src_valid~0_combout ),
	.src_valid1(\mm_interconnect_0|cmd_mux_010|src_valid~1_combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_010|src_data[46]~combout ),
	.out_data_buffer_65(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[65]~q ),
	.p1_wr_strobe(\epcs|the_niosII_epcs_sub|p1_wr_strobe~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_010|src_payload~2_combout ),
	.d_writedata_0(\cpu|cpu|d_writedata[0]~q ),
	.d_byteenable_0(\cpu|cpu|d_byteenable[0]~q ),
	.Equal9(\mm_interconnect_0|router|Equal9~0_combout ),
	.read_latency_shift_reg(\mm_interconnect_0|port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg~0_combout ),
	.d_writedata_1(\cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\cpu|cpu|d_writedata[7]~q ),
	.out_data_buffer_0(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[0]~q ),
	.out_data_toggle_flopped(\mm_interconnect_0|crosser_002|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\mm_interconnect_0|crosser_002|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.mem_used_12(\mm_interconnect_0|sys_pll_pll_slave_agent_rsp_fifo|mem_used[1]~q ),
	.wire_pfdena_reg_ena(\sys_pll|wire_pfdena_reg_ena~0_combout ),
	.out_data_buffer_651(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[65]~q ),
	.out_data_buffer_381(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_39(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[39]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.saved_grant_01(\mm_interconnect_0|cmd_mux_012|saved_grant[0]~q ),
	.d_byteenable_1(\cpu|cpu|d_byteenable[1]~q ),
	.use_reg(\mm_interconnect_0|sdram_s1_cmd_width_adapter|use_reg~q ),
	.saved_grant_11(\mm_interconnect_0|cmd_mux_012|saved_grant[1]~q ),
	.WideOr0(\mm_interconnect_0|sdram_s1_agent|WideOr0~2_combout ),
	.Equal0(\sdram|the_niosII_sdram_input_efifo_module|Equal0~0_combout ),
	.i_read(\cpu|cpu|i_read~q ),
	.F_pc_24(\cpu|cpu|F_pc[24]~q ),
	.F_pc_23(\cpu|cpu|F_pc[23]~q ),
	.F_pc_22(\cpu|cpu|F_pc[22]~q ),
	.F_pc_21(\cpu|cpu|F_pc[21]~q ),
	.F_pc_20(\cpu|cpu|F_pc[20]~q ),
	.F_pc_19(\cpu|cpu|F_pc[19]~q ),
	.F_pc_18(\cpu|cpu|F_pc[18]~q ),
	.F_pc_17(\cpu|cpu|F_pc[17]~q ),
	.F_pc_16(\cpu|cpu|F_pc[16]~q ),
	.F_pc_15(\cpu|cpu|F_pc[15]~q ),
	.F_pc_14(\cpu|cpu|F_pc[14]~q ),
	.F_pc_13(\cpu|cpu|F_pc[13]~q ),
	.F_pc_12(\cpu|cpu|F_pc[12]~q ),
	.F_pc_11(\cpu|cpu|F_pc[11]~q ),
	.F_pc_10(\cpu|cpu|F_pc[10]~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~0_combout ),
	.Equal4(\mm_interconnect_0|router|Equal4~1_combout ),
	.WideOr1(\mm_interconnect_0|cmd_mux_012|WideOr1~combout ),
	.m0_write1(\mm_interconnect_0|sdram_s1_agent|m0_write~2_combout ),
	.mem_used_7(\mm_interconnect_0|sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.src_data_66(\mm_interconnect_0|cmd_mux_012|src_data[66]~combout ),
	.F_pc_8(\cpu|cpu|F_pc[8]~q ),
	.out_data_28(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[28]~0_combout ),
	.src_valid2(\mm_interconnect_0|cmd_mux_012|src_valid~0_combout ),
	.src12_valid(\mm_interconnect_0|cmd_demux|src12_valid~0_combout ),
	.m0_write2(\mm_interconnect_0|sdram_s1_agent|m0_write~combout ),
	.out_data_42(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[42]~1_combout ),
	.F_pc_9(\cpu|cpu|F_pc[9]~q ),
	.out_data_29(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[29]~2_combout ),
	.out_data_31(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[31]~3_combout ),
	.out_data_30(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[30]~4_combout ),
	.out_data_33(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[33]~5_combout ),
	.out_data_32(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[32]~6_combout ),
	.out_data_35(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[35]~7_combout ),
	.out_data_34(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[34]~8_combout ),
	.out_data_37(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[37]~9_combout ),
	.out_data_36(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[36]~10_combout ),
	.out_data_39(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[39]~11_combout ),
	.out_data_38(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[38]~12_combout ),
	.out_data_41(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[41]~13_combout ),
	.out_data_40(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[40]~14_combout ),
	.out_data_19(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[19]~15_combout ),
	.F_pc_0(\cpu|cpu|F_pc[0]~q ),
	.out_data_20(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[20]~16_combout ),
	.F_pc_1(\cpu|cpu|F_pc[1]~q ),
	.out_data_21(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[21]~17_combout ),
	.F_pc_2(\cpu|cpu|F_pc[2]~q ),
	.out_data_22(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[22]~18_combout ),
	.F_pc_3(\cpu|cpu|F_pc[3]~q ),
	.out_data_23(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[23]~19_combout ),
	.F_pc_4(\cpu|cpu|F_pc[4]~q ),
	.out_data_24(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[24]~20_combout ),
	.F_pc_5(\cpu|cpu|F_pc[5]~q ),
	.out_data_25(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[25]~21_combout ),
	.F_pc_6(\cpu|cpu|F_pc[6]~q ),
	.out_data_26(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[26]~22_combout ),
	.F_pc_7(\cpu|cpu|F_pc[7]~q ),
	.out_data_27(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[27]~23_combout ),
	.always0(\adc_0|always0~1_combout ),
	.waitrequest(\adc_0|waitrequest~0_combout ),
	.mem_84_0(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][84]~q ),
	.mem_66_0(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][66]~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_01(\mm_interconnect_0|port_gpio_0_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_02(\mm_interconnect_0|sys_id_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_54_0(\mm_interconnect_0|sdram_s1_agent_rsp_fifo|mem[0][54]~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux_012|src0_valid~0_combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.mem_used_13(\mm_interconnect_0|timer_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|timer_0_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_11(\mm_interconnect_0|timer_0_s1_translator|wait_latency_counter[1]~q ),
	.read_latency_shift_reg1(\mm_interconnect_0|rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg~2_combout ),
	.write(\mm_interconnect_0|port_sw_avalon_parallel_port_slave_agent_rsp_fifo|write~2_combout ),
	.Equal12(\mm_interconnect_0|router|Equal12~1_combout ),
	.mem_used_14(\mm_interconnect_0|rs232_0_avalon_rs232_slave_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_02(\mm_interconnect_0|cmd_mux_009|saved_grant[0]~q ),
	.waitrequest1(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_15(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.cpu_data_master_waitrequest(\mm_interconnect_0|cpu_data_master_translator|av_waitrequest~1_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_010|src_payload~3_combout ),
	.src_data_661(\mm_interconnect_0|cmd_mux_010|src_data[66]~combout ),
	.av_begintransfer(\mm_interconnect_0|epcs_epcs_control_port_translator|av_begintransfer~0_combout ),
	.d_writedata_10(\cpu|cpu|d_writedata[10]~q ),
	.src_payload4(\mm_interconnect_0|cmd_mux_010|src_payload~4_combout ),
	.rst1(\jtag|niosII_jtag_alt_jtag_atlantic|rst1~q ),
	.out_data_buffer_66(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[66]~q ),
	.d_byteenable_2(\cpu|cpu|d_byteenable[2]~q ),
	.d_byteenable_3(\cpu|cpu|d_byteenable[3]~q ),
	.src1_valid(\mm_interconnect_0|rsp_demux_009|src1_valid~0_combout ),
	.read_accepted1(\mm_interconnect_0|cpu_instruction_master_translator|read_accepted~2_combout ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_012|src1_valid~0_combout ),
	.hbreak_enabled(\cpu|cpu|hbreak_enabled~q ),
	.read_latency_shift_reg2(\mm_interconnect_0|port_gpio_0_avalon_parallel_port_slave_translator|read_latency_shift_reg~0_combout ),
	.d_writedata_8(\cpu|cpu|d_writedata[8]~q ),
	.d_writedata_9(\cpu|cpu|d_writedata[9]~q ),
	.d_writedata_11(\cpu|cpu|d_writedata[11]~q ),
	.d_writedata_12(\cpu|cpu|d_writedata[12]~q ),
	.d_writedata_13(\cpu|cpu|d_writedata[13]~q ),
	.d_writedata_14(\cpu|cpu|d_writedata[14]~q ),
	.d_writedata_15(\cpu|cpu|d_writedata[15]~q ),
	.d_writedata_16(\cpu|cpu|d_writedata[16]~q ),
	.d_writedata_17(\cpu|cpu|d_writedata[17]~q ),
	.d_writedata_18(\cpu|cpu|d_writedata[18]~q ),
	.d_writedata_19(\cpu|cpu|d_writedata[19]~q ),
	.d_writedata_20(\cpu|cpu|d_writedata[20]~q ),
	.d_writedata_21(\cpu|cpu|d_writedata[21]~q ),
	.d_writedata_22(\cpu|cpu|d_writedata[22]~q ),
	.d_writedata_23(\cpu|cpu|d_writedata[23]~q ),
	.WideOr12(\mm_interconnect_0|cmd_mux_009|WideOr1~combout ),
	.write1(\mm_interconnect_0|port_key_avalon_parallel_port_slave_agent_rsp_fifo|write~0_combout ),
	.Equal121(\mm_interconnect_0|router|Equal12~2_combout ),
	.rf_source_valid(\mm_interconnect_0|cpu_debug_mem_slave_agent|rf_source_valid~0_combout ),
	.uav_write(\mm_interconnect_0|cpu_data_master_translator|uav_write~0_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_010|src_payload~5_combout ),
	.out_valid(\mm_interconnect_0|crosser_006|clock_xer|out_valid~combout ),
	.av_readdata_pre_0(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.out_data_buffer_01(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[0]~q ),
	.data_reg_0(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[0]~q ),
	.out_payload_0(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[0]~q ),
	.source_addr_1(\mm_interconnect_0|sdram_s1_agent|uncompressor|source_addr[1]~0_combout ),
	.F_iw_0(\cpu|cpu|F_iw[0]~5_combout ),
	.av_readdata_pre_1(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_1(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[1]~q ),
	.out_payload_1(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[1]~q ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~16_combout ),
	.av_readdata_pre_2(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.out_data_buffer_2(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[2]~q ),
	.data_reg_2(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[2]~q ),
	.out_payload_2(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[2]~q ),
	.F_iw_2(\cpu|cpu|F_iw[2]~10_combout ),
	.av_readdata_pre_3(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.out_data_buffer_3(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[3]~q ),
	.out_payload_3(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[3]~q ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~17_combout ),
	.av_readdata_pre_4(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.out_data_buffer_4(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[4]~q ),
	.out_payload_4(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[4]~q ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~18_combout ),
	.read_latency_shift_reg3(\mm_interconnect_0|rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg~1_combout ),
	.b_full(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.out_data_0(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[0]~24_combout ),
	.out_data_1(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[1]~25_combout ),
	.out_data_2(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[2]~26_combout ),
	.out_data_3(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[3]~27_combout ),
	.out_data_4(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[4]~28_combout ),
	.out_data_5(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[5]~29_combout ),
	.out_data_6(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[6]~30_combout ),
	.out_data_7(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[7]~31_combout ),
	.out_data_8(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[8]~32_combout ),
	.out_data_9(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[9]~33_combout ),
	.out_data_10(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[10]~34_combout ),
	.out_data_11(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[11]~35_combout ),
	.out_data_12(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[12]~36_combout ),
	.out_data_13(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[13]~37_combout ),
	.out_data_14(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[14]~38_combout ),
	.out_data_15(\mm_interconnect_0|sdram_s1_cmd_width_adapter|out_data[15]~39_combout ),
	.period_l_wr_strobe(\timer_0|period_l_wr_strobe~2_combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_009|src_data[46]~combout ),
	.out_data_toggle_flopped1(\mm_interconnect_0|crosser|clock_xer|out_data_toggle_flopped~q ),
	.av_readdata_pre_11(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.out_data_buffer_11(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[11]~q ),
	.out_payload_11(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[11]~q ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[11]~19_combout ),
	.av_readdata_pre_13(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.out_data_buffer_13(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[13]~q ),
	.out_payload_13(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[13]~q ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~20_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.out_data_buffer_16(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[16]~q ),
	.src_payload6(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.av_readdata_pre_12(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.out_data_buffer_12(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[12]~q ),
	.data_reg_12(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[12]~q ),
	.out_payload_12(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[12]~q ),
	.F_iw_12(\cpu|cpu|F_iw[12]~23_combout ),
	.av_readdata_pre_5(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.out_data_buffer_5(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[5]~q ),
	.out_payload_5(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[5]~q ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~21_combout ),
	.av_readdata_pre_14(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.out_data_buffer_14(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[14]~q ),
	.data_reg_14(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[14]~q ),
	.out_payload_14(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[14]~q ),
	.F_iw_14(\cpu|cpu|F_iw[14]~28_combout ),
	.av_readdata_pre_15(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.out_data_buffer_15(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[15]~q ),
	.out_payload_15(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[15]~q ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~22_combout ),
	.av_readdata_pre_10(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.out_data_buffer_10(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[10]~q ),
	.data_reg_10(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[10]~q ),
	.out_payload_10(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[10]~q ),
	.F_iw_10(\cpu|cpu|F_iw[10]~33_combout ),
	.av_readdata_pre_9(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.out_data_buffer_9(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[9]~q ),
	.data_reg_9(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[9]~q ),
	.out_payload_9(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[9]~q ),
	.F_iw_9(\cpu|cpu|F_iw[9]~36_combout ),
	.av_readdata_pre_8(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.out_data_buffer_8(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[8]~q ),
	.data_reg_8(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[8]~q ),
	.out_payload_8(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[8]~q ),
	.F_iw_8(\cpu|cpu|F_iw[8]~39_combout ),
	.av_readdata_pre_7(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.out_data_buffer_7(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[7]~q ),
	.data_reg_7(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[7]~q ),
	.out_payload_7(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[7]~q ),
	.F_iw_7(\cpu|cpu|F_iw[7]~42_combout ),
	.av_readdata_pre_6(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.out_data_buffer_6(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[6]~q ),
	.data_reg_6(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[6]~q ),
	.out_payload_6(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[6]~q ),
	.F_iw_6(\cpu|cpu|F_iw[6]~45_combout ),
	.av_readdata_pre_21(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.out_data_buffer_21(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[21]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.out_data_buffer_30(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[30]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.out_data_buffer_29(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[29]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.out_data_buffer_28(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[28]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.out_data_buffer_27(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[27]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.out_data_buffer_26(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[26]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.out_data_buffer_25(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[25]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.out_data_buffer_24(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[24]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.out_data_buffer_23(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[23]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.out_data_buffer_22(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[22]~q ),
	.av_readdata_pre_20(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.out_data_buffer_20(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[20]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.out_data_buffer_19(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[19]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.out_data_buffer_18(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.out_data_buffer_17(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[17]~q ),
	.src_payload7(\mm_interconnect_0|cmd_mux_010|src_payload~6_combout ),
	.readdata_02(\port_led|readdata[0]~q ),
	.readdata_03(\port_sw|readdata[0]~q ),
	.readdata_04(\port_key|readdata[0]~q ),
	.readdata_05(\port_gpio_0|readdata[0]~q ),
	.out_valid1(\mm_interconnect_0|crosser_005|clock_xer|out_valid~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~30_combout ),
	.readdata_06(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[0]~q ),
	.readdata_12(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[1]~q ),
	.readdata_2(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[2]~q ),
	.readdata_3(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[3]~q ),
	.readdata_13(\port_led|readdata[1]~q ),
	.readdata_14(\port_sw|readdata[1]~q ),
	.readdata_15(\port_key|readdata[1]~q ),
	.readdata_110(\port_gpio_0|readdata[1]~q ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[1]~38_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~39_combout ),
	.readdata_24(\port_led|readdata[2]~q ),
	.readdata_25(\port_gpio_0|readdata[2]~q ),
	.readdata_26(\port_sw|readdata[2]~q ),
	.readdata_27(\rs232_1|readdata[2]~q ),
	.readdata_28(\rs232_0|readdata[2]~q ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[2]~45_combout ),
	.readdata_31(\port_led|readdata[3]~q ),
	.readdata_32(\port_gpio_0|readdata[3]~q ),
	.readdata_33(\port_sw|readdata[3]~q ),
	.readdata_34(\rs232_1|readdata[3]~q ),
	.readdata_35(\rs232_0|readdata[3]~q ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[3]~52_combout ),
	.readdata_41(\port_led|readdata[4]~q ),
	.readdata_42(\rs232_0|readdata[4]~q ),
	.readdata_43(\port_gpio_0|readdata[4]~q ),
	.readdata_44(\rs232_1|readdata[4]~q ),
	.av_readdata_pre_301(\mm_interconnect_0|sys_id_control_slave_translator|av_readdata_pre[30]~q ),
	.src_data_41(\mm_interconnect_0|rsp_mux|src_data[4]~58_combout ),
	.readdata_5(\port_led|readdata[5]~q ),
	.readdata_51(\rs232_0|readdata[5]~q ),
	.readdata_52(\port_gpio_0|readdata[5]~q ),
	.readdata_53(\rs232_1|readdata[5]~q ),
	.src_data_51(\mm_interconnect_0|rsp_mux|src_data[5]~64_combout ),
	.readdata_6(\port_led|readdata[6]~q ),
	.readdata_61(\rs232_0|readdata[6]~q ),
	.readdata_62(\port_gpio_0|readdata[6]~q ),
	.readdata_63(\rs232_1|readdata[6]~q ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~70_combout ),
	.readdata_7(\port_led|readdata[7]~q ),
	.readdata_71(\rs232_0|readdata[7]~q ),
	.readdata_72(\port_gpio_0|readdata[7]~q ),
	.readdata_73(\rs232_1|readdata[7]~q ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~76_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_009|src_payload~0_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_009|src_payload~1_combout ),
	.src_data_381(\mm_interconnect_0|cmd_mux_009|src_data[38]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux_009|src_data[39]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_009|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_009|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_009|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_009|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_009|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_009|src_data[45]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_009|src_data[32]~combout ),
	.b_non_empty(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_5(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag|the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.dreg_01(\mm_interconnect_0|crosser|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.av_waitrequest(\jtag|av_waitrequest~q ),
	.mem_used_16(\mm_interconnect_0|jtag_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.out_data_buffer_661(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[66]~q ),
	.out_data_buffer_382(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_71(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[7]~q ),
	.za_valid(\sdram|za_valid~q ),
	.readdata_111(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[11]~q ),
	.readdata_131(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[13]~q ),
	.readdata_162(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[16]~q ),
	.readdata_121(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[12]~q ),
	.readdata_54(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[5]~q ),
	.readdata_141(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[14]~q ),
	.readdata_151(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[15]~q ),
	.readdata_10(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[10]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.out_data_buffer_31(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[31]~q ),
	.readdata_9(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[9]~q ),
	.readdata_8(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[8]~q ),
	.readdata_74(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[7]~q ),
	.readdata_64(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[6]~q ),
	.out_data_buffer_261(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[26]~q ),
	.readdata_212(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[21]~q ),
	.readdata_30(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[30]~q ),
	.out_data_buffer_251(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[25]~q ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~5_combout ),
	.readdata_29(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[29]~q ),
	.out_data_buffer_241(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[24]~q ),
	.readdata_281(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[28]~q ),
	.readdata_232(\port_gpio_0|readdata[23]~q ),
	.src_payload11(\mm_interconnect_0|rsp_mux|src_payload~9_combout ),
	.readdata_271(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[27]~q ),
	.readdata_222(\port_gpio_0|readdata[22]~q ),
	.src_payload12(\mm_interconnect_0|rsp_mux|src_payload~14_combout ),
	.readdata_261(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[26]~q ),
	.readdata_213(\port_gpio_0|readdata[21]~q ),
	.src_payload13(\mm_interconnect_0|rsp_mux|src_payload~19_combout ),
	.readdata_251(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[25]~q ),
	.readdata_202(\port_gpio_0|readdata[20]~q ),
	.src_payload14(\mm_interconnect_0|rsp_mux|src_payload~24_combout ),
	.readdata_241(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[24]~q ),
	.readdata_192(\port_gpio_0|readdata[19]~q ),
	.src_payload15(\mm_interconnect_0|rsp_mux|src_payload~29_combout ),
	.readdata_233(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[23]~q ),
	.readdata_182(\port_gpio_0|readdata[18]~q ),
	.src_payload16(\mm_interconnect_0|rsp_mux|src_payload~34_combout ),
	.readdata_223(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[22]~q ),
	.readdata_172(\port_gpio_0|readdata[17]~q ),
	.src_payload17(\mm_interconnect_0|rsp_mux|src_payload~39_combout ),
	.readdata_163(\port_gpio_0|readdata[16]~q ),
	.src_payload18(\mm_interconnect_0|rsp_mux|src_payload~44_combout ),
	.readdata_203(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[20]~q ),
	.readdata_152(\port_gpio_0|readdata[15]~q ),
	.readdata_153(\rs232_1|readdata[15]~q ),
	.readdata_154(\rs232_0|readdata[15]~q ),
	.src_data_151(\mm_interconnect_0|rsp_mux|src_data[15]~82_combout ),
	.readdata_193(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[19]~q ),
	.readdata_142(\port_gpio_0|readdata[14]~q ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~85_combout ),
	.readdata_183(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[18]~q ),
	.readdata_132(\port_gpio_0|readdata[13]~q ),
	.src_data_131(\mm_interconnect_0|rsp_mux|src_data[13]~89_combout ),
	.readdata_173(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[17]~q ),
	.readdata_122(\port_gpio_0|readdata[12]~q ),
	.src_data_121(\mm_interconnect_0|rsp_mux|src_data[12]~92_combout ),
	.readdata_112(\port_gpio_0|readdata[11]~q ),
	.src_data_111(\mm_interconnect_0|rsp_mux|src_data[11]~96_combout ),
	.readdata_101(\port_gpio_0|readdata[10]~q ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~101_combout ),
	.readdata_91(\port_gpio_0|readdata[9]~q ),
	.readdata_92(\rs232_1|readdata[9]~q ),
	.readdata_93(\rs232_0|readdata[9]~q ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~107_combout ),
	.readdata_81(\port_gpio_0|readdata[8]~q ),
	.readdata_82(\rs232_1|readdata[8]~q ),
	.readdata_83(\rs232_0|readdata[8]~q ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~113_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_010|src_payload~7_combout ),
	.av_readdata_pre_01(\mm_interconnect_0|adc_0_adc_slave_translator|av_readdata_pre[0]~0_combout ),
	.readdata_07(\adc_0|readdata[0]~4_combout ),
	.readdata_08(\timer_0|readdata[0]~q ),
	.readdata_113(\adc_0|readdata[1]~9_combout ),
	.readdata_114(\timer_0|readdata[1]~q ),
	.readdata_210(\adc_0|readdata[2]~14_combout ),
	.readdata_214(\timer_0|readdata[2]~q ),
	.readdata_36(\adc_0|readdata[3]~19_combout ),
	.readdata_37(\timer_0|readdata[3]~q ),
	.readdata_45(\adc_0|readdata[4]~24_combout ),
	.readdata_46(\timer_0|readdata[4]~q ),
	.readdata_55(\adc_0|readdata[5]~29_combout ),
	.readdata_56(\timer_0|readdata[5]~q ),
	.readdata_65(\adc_0|readdata[6]~34_combout ),
	.readdata_66(\timer_0|readdata[6]~q ),
	.readdata_75(\adc_0|readdata[7]~39_combout ),
	.readdata_76(\timer_0|readdata[7]~q ),
	.src_payload20(\mm_interconnect_0|cmd_mux_009|src_payload~2_combout ),
	.out_data_buffer_652(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[65]~q ),
	.out_data_buffer_02(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[0]~q ),
	.b_full1(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_21(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_11(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_51(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_41(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_31(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_01(\jtag|the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.out_data_buffer_271(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_281(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[28]~q ),
	.out_data_buffer_291(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_301(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[30]~q ),
	.out_data_buffer_311(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[31]~q ),
	.readdata_311(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[31]~q ),
	.readdata_155(\adc_0|readdata[15]~40_combout ),
	.readdata_156(\timer_0|readdata[15]~q ),
	.readdata_143(\timer_0|readdata[14]~q ),
	.readdata_133(\timer_0|readdata[13]~q ),
	.readdata_123(\timer_0|readdata[12]~q ),
	.readdata_115(\adc_0|readdata[11]~45_combout ),
	.readdata_116(\timer_0|readdata[11]~q ),
	.readdata_102(\timer_0|readdata[10]~q ),
	.readdata_103(\adc_0|readdata[10]~50_combout ),
	.readdata_94(\adc_0|readdata[9]~55_combout ),
	.readdata_95(\timer_0|readdata[9]~q ),
	.readdata_84(\adc_0|readdata[8]~60_combout ),
	.readdata_85(\timer_0|readdata[8]~q ),
	.src_payload21(\mm_interconnect_0|cmd_mux_010|src_payload~8_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_009|src_payload~3_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_009|src_payload~4_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_009|src_payload~5_combout ),
	.readdata_09(\epcs|readdata[0]~0_combout ),
	.za_data_0(\sdram|za_data[0]~q ),
	.readdata_117(\epcs|readdata[1]~1_combout ),
	.za_data_1(\sdram|za_data[1]~q ),
	.readdata_215(\epcs|readdata[2]~2_combout ),
	.za_data_2(\sdram|za_data[2]~q ),
	.readdata_38(\epcs|readdata[3]~3_combout ),
	.za_data_3(\sdram|za_data[3]~q ),
	.readdata_47(\epcs|readdata[4]~4_combout ),
	.za_data_4(\sdram|za_data[4]~q ),
	.out_data_buffer_110(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[1]~q ),
	.readdata_118(\epcs|readdata[11]~5_combout ),
	.za_data_11(\sdram|za_data[11]~q ),
	.readdata_134(\epcs|readdata[13]~6_combout ),
	.za_data_13(\sdram|za_data[13]~q ),
	.readdata_164(\epcs|readdata[16]~7_combout ),
	.readdata_124(\epcs|readdata[12]~8_combout ),
	.za_data_12(\sdram|za_data[12]~q ),
	.readdata_57(\epcs|readdata[5]~9_combout ),
	.za_data_5(\sdram|za_data[5]~q ),
	.readdata_144(\epcs|readdata[14]~10_combout ),
	.za_data_14(\sdram|za_data[14]~q ),
	.readdata_157(\epcs|readdata[15]~11_combout ),
	.za_data_15(\sdram|za_data[15]~q ),
	.readdata_104(\epcs|readdata[10]~12_combout ),
	.za_data_10(\sdram|za_data[10]~q ),
	.readdata_96(\epcs|readdata[9]~13_combout ),
	.za_data_9(\sdram|za_data[9]~q ),
	.readdata_86(\epcs|readdata[8]~14_combout ),
	.za_data_8(\sdram|za_data[8]~q ),
	.readdata_77(\epcs|readdata[7]~15_combout ),
	.za_data_7(\sdram|za_data[7]~q ),
	.readdata_67(\epcs|readdata[6]~16_combout ),
	.za_data_6(\sdram|za_data[6]~q ),
	.readdata_216(\epcs|readdata[21]~17_combout ),
	.readdata_301(\epcs|readdata[30]~18_combout ),
	.readdata_291(\epcs|readdata[29]~19_combout ),
	.readdata_282(\epcs|readdata[28]~20_combout ),
	.readdata_272(\epcs|readdata[27]~21_combout ),
	.readdata_262(\epcs|readdata[26]~22_combout ),
	.readdata_252(\epcs|readdata[25]~23_combout ),
	.readdata_242(\epcs|readdata[24]~24_combout ),
	.readdata_234(\epcs|readdata[23]~25_combout ),
	.readdata_224(\epcs|readdata[22]~26_combout ),
	.readdata_204(\epcs|readdata[20]~27_combout ),
	.readdata_194(\epcs|readdata[19]~28_combout ),
	.readdata_184(\epcs|readdata[18]~29_combout ),
	.readdata_174(\epcs|readdata[17]~30_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_010|src_payload~9_combout ),
	.read_0(\jtag|read_0~q ),
	.av_readdata_0(\jtag|av_readdata[0]~0_combout ),
	.readdata_010(\sys_pll|readdata[0]~1_combout ),
	.av_readdata_9(\jtag|av_readdata[9]~combout ),
	.src_data_412(\mm_interconnect_0|cmd_mux_010|src_data[41]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_010|src_data[42]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_010|src_data[43]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_010|src_data[44]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_010|src_data[45]~combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_010|src_payload~10_combout ),
	.av_readdata_1(\jtag|av_readdata[1]~1_combout ),
	.readdata_119(\sys_pll|readdata[1]~2_combout ),
	.av_readdata_2(\jtag|av_readdata[2]~2_combout ),
	.av_readdata_3(\jtag|av_readdata[3]~3_combout ),
	.av_readdata_4(\jtag|av_readdata[4]~4_combout ),
	.av_readdata_5(\jtag|av_readdata[5]~5_combout ),
	.av_readdata_6(\jtag|av_readdata[6]~6_combout ),
	.av_readdata_7(\jtag|av_readdata[7]~7_combout ),
	.out_data_buffer_210(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[2]~q ),
	.src_payload27(\mm_interconnect_0|cmd_mux_009|src_payload~6_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_009|src_data[33]~combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_009|src_payload~7_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_009|src_payload~8_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_009|src_data[34]~combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_009|src_payload~9_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_009|src_payload~10_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_009|src_payload~11_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_009|src_payload~12_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_009|src_payload~13_combout ),
	.readdata_312(\epcs|readdata[31]~31_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_009|src_payload~14_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_009|src_payload~15_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_009|src_payload~16_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_009|src_payload~17_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_009|src_payload~18_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_009|src_payload~19_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_009|src_data[35]~combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_009|src_payload~20_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_009|src_payload~21_combout ),
	.src_payload43(\mm_interconnect_0|cmd_mux_009|src_payload~22_combout ),
	.src_payload44(\mm_interconnect_0|cmd_mux_009|src_payload~23_combout ),
	.src_payload45(\mm_interconnect_0|cmd_mux_009|src_payload~24_combout ),
	.src_payload46(\mm_interconnect_0|cmd_mux_009|src_payload~25_combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_009|src_payload~26_combout ),
	.src_payload48(\mm_interconnect_0|cmd_mux_009|src_payload~27_combout ),
	.src_payload49(\mm_interconnect_0|cmd_mux_009|src_payload~28_combout ),
	.rvalid(\jtag|rvalid~q ),
	.src_payload50(\mm_interconnect_0|cmd_mux_009|src_payload~29_combout ),
	.woverflow(\jtag|woverflow~q ),
	.src_payload51(\mm_interconnect_0|cmd_mux_009|src_payload~30_combout ),
	.src_payload52(\mm_interconnect_0|cmd_mux_009|src_payload~31_combout ),
	.ac(\jtag|ac~q ),
	.av_readdata_8(\jtag|av_readdata[8]~8_combout ),
	.out_data_buffer_111(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_32(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[3]~q ),
	.src_payload53(\mm_interconnect_0|cmd_mux_010|src_payload~11_combout ),
	.src_payload54(\mm_interconnect_0|cmd_mux_010|src_payload~12_combout ),
	.src_payload55(\mm_interconnect_0|cmd_mux_010|src_payload~13_combout ),
	.src_payload56(\mm_interconnect_0|cmd_mux_010|src_payload~14_combout ),
	.src_payload57(\mm_interconnect_0|cmd_mux_010|src_payload~15_combout ),
	.src_payload58(\mm_interconnect_0|cmd_mux_009|src_payload~32_combout ),
	.src_payload59(\mm_interconnect_0|cmd_mux_010|src_payload~16_combout ),
	.src_payload60(\mm_interconnect_0|cmd_mux_010|src_payload~17_combout ),
	.out_data_buffer_101(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_41(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_51(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_61(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[6]~q ),
	.write2(\mm_interconnect_0|port_sw_avalon_parallel_port_slave_agent_rsp_fifo|write~3_combout ),
	.clk_clk(\clk_clk~input_o ));

niosII_niosII_timer_0 timer_0(
	.clk(\sys_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_4(\cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.hold_waitrequest(\mm_interconnect_0|cpu_data_master_agent|hold_waitrequest~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|cpu_data_master_translator|write_accepted~q ),
	.read_mux_out(\timer_0|read_mux_out~0_combout ),
	.writedata({\cpu|cpu|d_writedata[15]~q ,\cpu|cpu|d_writedata[14]~q ,\cpu|cpu|d_writedata[13]~q ,\cpu|cpu|d_writedata[12]~q ,\cpu|cpu|d_writedata[11]~q ,\cpu|cpu|d_writedata[10]~q ,\cpu|cpu|d_writedata[9]~q ,\cpu|cpu|d_writedata[8]~q ,\cpu|cpu|d_writedata[7]~q ,
\cpu|cpu|d_writedata[6]~q ,\cpu|cpu|d_writedata[5]~q ,\cpu|cpu|d_writedata[4]~q ,\cpu|cpu|d_writedata[3]~q ,\cpu|cpu|d_writedata[2]~q ,\cpu|cpu|d_writedata[1]~q ,\cpu|cpu|d_writedata[0]~q }),
	.Equal6(\timer_0|Equal6~0_combout ),
	.Equal4(\mm_interconnect_0|router|Equal4~1_combout ),
	.mem_used_1(\mm_interconnect_0|timer_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|timer_0_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|timer_0_s1_translator|wait_latency_counter[1]~q ),
	.Equal61(\timer_0|Equal6~1_combout ),
	.uav_write(\mm_interconnect_0|cpu_data_master_translator|uav_write~0_combout ),
	.period_l_wr_strobe1(\timer_0|period_l_wr_strobe~2_combout ),
	.timeout_occurred1(\timer_0|timeout_occurred~q ),
	.control_register_0(\timer_0|control_register[0]~q ),
	.readdata_0(\timer_0|readdata[0]~q ),
	.readdata_1(\timer_0|readdata[1]~q ),
	.readdata_2(\timer_0|readdata[2]~q ),
	.readdata_3(\timer_0|readdata[3]~q ),
	.readdata_4(\timer_0|readdata[4]~q ),
	.readdata_5(\timer_0|readdata[5]~q ),
	.readdata_6(\timer_0|readdata[6]~q ),
	.readdata_7(\timer_0|readdata[7]~q ),
	.readdata_15(\timer_0|readdata[15]~q ),
	.readdata_14(\timer_0|readdata[14]~q ),
	.readdata_13(\timer_0|readdata[13]~q ),
	.readdata_12(\timer_0|readdata[12]~q ),
	.readdata_11(\timer_0|readdata[11]~q ),
	.readdata_10(\timer_0|readdata[10]~q ),
	.readdata_9(\timer_0|readdata[9]~q ),
	.readdata_8(\timer_0|readdata[8]~q ));

niosII_niosII_sys_pll sys_pll(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.wire_pll7_clk_1(\sys_pll|sd1|wire_pll7_clk[1] ),
	.out_data_buffer_0(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[0]~q ),
	.out_data_toggle_flopped(\mm_interconnect_0|crosser_002|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\mm_interconnect_0|crosser_002|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.mem_used_1(\mm_interconnect_0|sys_pll_pll_slave_agent_rsp_fifo|mem_used[1]~q ),
	.wire_pfdena_reg_ena(\sys_pll|wire_pfdena_reg_ena~0_combout ),
	.out_data_buffer_65(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[65]~q ),
	.out_data_buffer_38(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_39(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[39]~q ),
	.reset(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.out_data_buffer_66(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[66]~q ),
	.readdata_0(\sys_pll|readdata[0]~1_combout ),
	.readdata_1(\sys_pll|readdata[1]~2_combout ),
	.out_data_buffer_1(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[1]~q ),
	.clk_clk(\clk_clk~input_o ));

niosII_altera_reset_controller rst_controller(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.reset_reset_n(\reset_reset_n~input_o ));

niosII_altera_irq_clock_crosser_1 irq_synchronizer_001(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.dreg_1(\irq_synchronizer_001|sync|sync[0].u|dreg[1]~q ),
	.irq_reg(\epcs|the_niosII_epcs_sub|irq_reg~q ));

niosII_altera_irq_clock_crosser irq_synchronizer(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.dreg_1(\irq_synchronizer|sync|sync[0].u|dreg[1]~q ),
	.av_irq(\jtag|av_irq~combout ));

niosII_altera_reset_controller_2 rst_controller_002(
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

niosII_altera_reset_controller_1 rst_controller_001(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.r_sync_rst1(\rst_controller_001|r_sync_rst~q ),
	.resetrequest(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_oci_debug|resetrequest~q ),
	.r_early_rst1(\rst_controller_001|r_early_rst~q ),
	.reset_reset_n(\reset_reset_n~input_o ));

niosII_niosII_cpu cpu(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.sr_0(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.W_alu_result_6(\cpu|cpu|W_alu_result[6]~q ),
	.W_alu_result_26(\cpu|cpu|W_alu_result[26]~q ),
	.W_alu_result_25(\cpu|cpu|W_alu_result[25]~q ),
	.W_alu_result_24(\cpu|cpu|W_alu_result[24]~q ),
	.W_alu_result_23(\cpu|cpu|W_alu_result[23]~q ),
	.W_alu_result_22(\cpu|cpu|W_alu_result[22]~q ),
	.W_alu_result_21(\cpu|cpu|W_alu_result[21]~q ),
	.W_alu_result_20(\cpu|cpu|W_alu_result[20]~q ),
	.W_alu_result_19(\cpu|cpu|W_alu_result[19]~q ),
	.W_alu_result_18(\cpu|cpu|W_alu_result[18]~q ),
	.W_alu_result_17(\cpu|cpu|W_alu_result[17]~q ),
	.W_alu_result_16(\cpu|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\cpu|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\cpu|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\cpu|cpu|W_alu_result[13]~q ),
	.W_alu_result_12(\cpu|cpu|W_alu_result[12]~q ),
	.W_alu_result_11(\cpu|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\cpu|cpu|W_alu_result[10]~q ),
	.W_alu_result_5(\cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_7(\cpu|cpu|W_alu_result[7]~q ),
	.W_alu_result_9(\cpu|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\cpu|cpu|W_alu_result[8]~q ),
	.W_alu_result_4(\cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.d_writedata_24(\cpu|cpu|d_writedata[24]~q ),
	.d_writedata_25(\cpu|cpu|d_writedata[25]~q ),
	.d_writedata_26(\cpu|cpu|d_writedata[26]~q ),
	.d_writedata_27(\cpu|cpu|d_writedata[27]~q ),
	.d_writedata_28(\cpu|cpu|d_writedata[28]~q ),
	.d_writedata_29(\cpu|cpu|d_writedata[29]~q ),
	.d_writedata_30(\cpu|cpu|d_writedata[30]~q ),
	.d_writedata_31(\cpu|cpu|d_writedata[31]~q ),
	.irq(\rs232_1|irq~q ),
	.irq1(\rs232_0|irq~q ),
	.readdata_4(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[4]~q ),
	.ir_out_0(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|ir_out[0]~q ),
	.ir_out_1(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|ir_out[1]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_read(\cpu|cpu|d_read~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.d_writedata_0(\cpu|cpu|d_writedata[0]~q ),
	.d_byteenable_0(\cpu|cpu|d_byteenable[0]~q ),
	.d_writedata_1(\cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\cpu|cpu|d_writedata[7]~q ),
	.d_byteenable_1(\cpu|cpu|d_byteenable[1]~q ),
	.i_read(\cpu|cpu|i_read~q ),
	.F_pc_24(\cpu|cpu|F_pc[24]~q ),
	.F_pc_23(\cpu|cpu|F_pc[23]~q ),
	.F_pc_22(\cpu|cpu|F_pc[22]~q ),
	.F_pc_21(\cpu|cpu|F_pc[21]~q ),
	.F_pc_20(\cpu|cpu|F_pc[20]~q ),
	.F_pc_19(\cpu|cpu|F_pc[19]~q ),
	.F_pc_18(\cpu|cpu|F_pc[18]~q ),
	.F_pc_17(\cpu|cpu|F_pc[17]~q ),
	.F_pc_16(\cpu|cpu|F_pc[16]~q ),
	.F_pc_15(\cpu|cpu|F_pc[15]~q ),
	.F_pc_14(\cpu|cpu|F_pc[14]~q ),
	.F_pc_13(\cpu|cpu|F_pc[13]~q ),
	.F_pc_12(\cpu|cpu|F_pc[12]~q ),
	.F_pc_11(\cpu|cpu|F_pc[11]~q ),
	.F_pc_10(\cpu|cpu|F_pc[10]~q ),
	.F_pc_8(\cpu|cpu|F_pc[8]~q ),
	.F_pc_9(\cpu|cpu|F_pc[9]~q ),
	.F_pc_0(\cpu|cpu|F_pc[0]~q ),
	.F_pc_1(\cpu|cpu|F_pc[1]~q ),
	.F_pc_2(\cpu|cpu|F_pc[2]~q ),
	.F_pc_3(\cpu|cpu|F_pc[3]~q ),
	.F_pc_4(\cpu|cpu|F_pc[4]~q ),
	.F_pc_5(\cpu|cpu|F_pc[5]~q ),
	.F_pc_6(\cpu|cpu|F_pc[6]~q ),
	.F_pc_7(\cpu|cpu|F_pc[7]~q ),
	.mem_84_0(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][84]~q ),
	.mem_66_0(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][66]~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_01(\mm_interconnect_0|port_gpio_0_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_02(\mm_interconnect_0|sys_id_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_54_0(\mm_interconnect_0|sdram_s1_agent_rsp_fifo|mem[0][54]~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux_012|src0_valid~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_009|saved_grant[0]~q ),
	.debug_mem_slave_waitrequest(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(\mm_interconnect_0|cpu_data_master_translator|av_waitrequest~1_combout ),
	.d_writedata_10(\cpu|cpu|d_writedata[10]~q ),
	.d_byteenable_2(\cpu|cpu|d_byteenable[2]~q ),
	.d_byteenable_3(\cpu|cpu|d_byteenable[3]~q ),
	.src1_valid(\mm_interconnect_0|rsp_demux_009|src1_valid~0_combout ),
	.read_accepted(\mm_interconnect_0|cpu_instruction_master_translator|read_accepted~2_combout ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_012|src1_valid~0_combout ),
	.hbreak_enabled(\cpu|cpu|hbreak_enabled~q ),
	.d_writedata_8(\cpu|cpu|d_writedata[8]~q ),
	.d_writedata_9(\cpu|cpu|d_writedata[9]~q ),
	.d_writedata_11(\cpu|cpu|d_writedata[11]~q ),
	.d_writedata_12(\cpu|cpu|d_writedata[12]~q ),
	.d_writedata_13(\cpu|cpu|d_writedata[13]~q ),
	.d_writedata_14(\cpu|cpu|d_writedata[14]~q ),
	.d_writedata_15(\cpu|cpu|d_writedata[15]~q ),
	.d_writedata_16(\cpu|cpu|d_writedata[16]~q ),
	.d_writedata_17(\cpu|cpu|d_writedata[17]~q ),
	.d_writedata_18(\cpu|cpu|d_writedata[18]~q ),
	.d_writedata_19(\cpu|cpu|d_writedata[19]~q ),
	.d_writedata_20(\cpu|cpu|d_writedata[20]~q ),
	.d_writedata_21(\cpu|cpu|d_writedata[21]~q ),
	.d_writedata_22(\cpu|cpu|d_writedata[22]~q ),
	.d_writedata_23(\cpu|cpu|d_writedata[23]~q ),
	.WideOr11(\mm_interconnect_0|cmd_mux_009|WideOr1~combout ),
	.rf_source_valid(\mm_interconnect_0|cpu_debug_mem_slave_agent|rf_source_valid~0_combout ),
	.uav_write(\mm_interconnect_0|cpu_data_master_translator|uav_write~0_combout ),
	.out_valid(\mm_interconnect_0|crosser_006|clock_xer|out_valid~combout ),
	.av_readdata_pre_0(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.out_data_buffer_0(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[0]~q ),
	.data_reg_0(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[0]~q ),
	.out_payload_0(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[0]~q ),
	.source_addr_1(\mm_interconnect_0|sdram_s1_agent|uncompressor|source_addr[1]~0_combout ),
	.F_iw_0(\cpu|cpu|F_iw[0]~5_combout ),
	.av_readdata_pre_1(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_1(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[1]~q ),
	.out_payload_1(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[1]~q ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~16_combout ),
	.av_readdata_pre_2(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.out_data_buffer_2(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[2]~q ),
	.data_reg_2(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[2]~q ),
	.out_payload_2(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[2]~q ),
	.F_iw_2(\cpu|cpu|F_iw[2]~10_combout ),
	.av_readdata_pre_3(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.out_data_buffer_3(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[3]~q ),
	.out_payload_3(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[3]~q ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~17_combout ),
	.av_readdata_pre_4(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.out_data_buffer_4(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[4]~q ),
	.out_payload_4(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[4]~q ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~18_combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_009|src_data[46]~combout ),
	.av_readdata_pre_11(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.out_data_buffer_11(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[11]~q ),
	.out_payload_11(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[11]~q ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[11]~19_combout ),
	.av_readdata_pre_13(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.out_data_buffer_13(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[13]~q ),
	.out_payload_13(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[13]~q ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~20_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.out_data_buffer_16(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[16]~q ),
	.src_payload(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.av_readdata_pre_12(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.out_data_buffer_12(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[12]~q ),
	.data_reg_12(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[12]~q ),
	.out_payload_12(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[12]~q ),
	.F_iw_12(\cpu|cpu|F_iw[12]~23_combout ),
	.av_readdata_pre_5(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.out_data_buffer_5(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[5]~q ),
	.out_payload_5(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[5]~q ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~21_combout ),
	.av_readdata_pre_14(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.out_data_buffer_14(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[14]~q ),
	.data_reg_14(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[14]~q ),
	.out_payload_14(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[14]~q ),
	.F_iw_14(\cpu|cpu|F_iw[14]~28_combout ),
	.av_readdata_pre_15(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.out_data_buffer_15(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[15]~q ),
	.out_payload_15(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[15]~q ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~22_combout ),
	.av_readdata_pre_10(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.out_data_buffer_10(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[10]~q ),
	.data_reg_10(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[10]~q ),
	.out_payload_10(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[10]~q ),
	.F_iw_10(\cpu|cpu|F_iw[10]~33_combout ),
	.av_readdata_pre_9(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.out_data_buffer_9(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[9]~q ),
	.data_reg_9(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[9]~q ),
	.out_payload_9(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[9]~q ),
	.F_iw_9(\cpu|cpu|F_iw[9]~36_combout ),
	.av_readdata_pre_8(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.out_data_buffer_8(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[8]~q ),
	.data_reg_8(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[8]~q ),
	.out_payload_8(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[8]~q ),
	.F_iw_8(\cpu|cpu|F_iw[8]~39_combout ),
	.av_readdata_pre_7(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.out_data_buffer_7(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[7]~q ),
	.data_reg_7(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[7]~q ),
	.out_payload_7(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[7]~q ),
	.F_iw_7(\cpu|cpu|F_iw[7]~42_combout ),
	.av_readdata_pre_6(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.out_data_buffer_6(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[6]~q ),
	.data_reg_6(\mm_interconnect_0|sdram_s1_rsp_width_adapter|data_reg[6]~q ),
	.out_payload_6(\mm_interconnect_0|sdram_s1_agent_rdata_fifo|out_payload[6]~q ),
	.F_iw_6(\cpu|cpu|F_iw[6]~45_combout ),
	.av_readdata_pre_21(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.out_data_buffer_21(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[21]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.out_data_buffer_30(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[30]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.out_data_buffer_29(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[29]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.out_data_buffer_28(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[28]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.out_data_buffer_27(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[27]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.out_data_buffer_26(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[26]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.out_data_buffer_25(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[25]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.out_data_buffer_24(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[24]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.out_data_buffer_23(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[23]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.out_data_buffer_22(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[22]~q ),
	.av_readdata_pre_20(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.out_data_buffer_20(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[20]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.out_data_buffer_19(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[19]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.out_data_buffer_18(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.out_data_buffer_17(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[17]~q ),
	.out_valid1(\mm_interconnect_0|crosser_005|clock_xer|out_valid~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~30_combout ),
	.dreg_1(\irq_synchronizer_001|sync|sync[0].u|dreg[1]~q ),
	.timeout_occurred(\timer_0|timeout_occurred~q ),
	.control_register_0(\timer_0|control_register[0]~q ),
	.dreg_11(\irq_synchronizer|sync|sync[0].u|dreg[1]~q ),
	.readdata_0(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[0]~q ),
	.readdata_1(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[1]~q ),
	.readdata_2(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[2]~q ),
	.readdata_3(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[3]~q ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[1]~38_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~39_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[2]~45_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[3]~52_combout ),
	.av_readdata_pre_301(\mm_interconnect_0|sys_id_control_slave_translator|av_readdata_pre[30]~q ),
	.src_data_41(\mm_interconnect_0|rsp_mux|src_data[4]~58_combout ),
	.src_data_51(\mm_interconnect_0|rsp_mux|src_data[5]~64_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~70_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~76_combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_009|src_payload~0_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_009|src_payload~1_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_009|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_009|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_009|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_009|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_009|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_009|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_009|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_009|src_data[45]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_009|src_data[32]~combout ),
	.readdata_11(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[11]~q ),
	.readdata_13(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[13]~q ),
	.readdata_16(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[16]~q ),
	.readdata_12(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[12]~q ),
	.readdata_5(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[5]~q ),
	.readdata_14(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[14]~q ),
	.readdata_15(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[15]~q ),
	.readdata_10(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[10]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.out_data_buffer_31(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[31]~q ),
	.readdata_9(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[9]~q ),
	.readdata_8(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[8]~q ),
	.readdata_7(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[7]~q ),
	.readdata_6(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[6]~q ),
	.readdata_26(\port_gpio_0|readdata[26]~q ),
	.out_data_buffer_261(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[26]~q ),
	.readdata_21(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[21]~q ),
	.readdata_30(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[30]~q ),
	.readdata_25(\port_gpio_0|readdata[25]~q ),
	.out_data_buffer_251(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[25]~q ),
	.src_payload3(\mm_interconnect_0|rsp_mux|src_payload~5_combout ),
	.readdata_29(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[29]~q ),
	.readdata_24(\port_gpio_0|readdata[24]~q ),
	.out_data_buffer_241(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[24]~q ),
	.readdata_28(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[28]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~9_combout ),
	.readdata_27(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[27]~q ),
	.src_payload5(\mm_interconnect_0|rsp_mux|src_payload~14_combout ),
	.readdata_261(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[26]~q ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~19_combout ),
	.readdata_251(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[25]~q ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~24_combout ),
	.readdata_241(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[24]~q ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~29_combout ),
	.readdata_23(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[23]~q ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~34_combout ),
	.readdata_22(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[22]~q ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~39_combout ),
	.src_payload11(\mm_interconnect_0|rsp_mux|src_payload~44_combout ),
	.readdata_20(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[20]~q ),
	.src_data_151(\mm_interconnect_0|rsp_mux|src_data[15]~82_combout ),
	.readdata_19(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[19]~q ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~85_combout ),
	.readdata_18(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[18]~q ),
	.src_data_131(\mm_interconnect_0|rsp_mux|src_data[13]~89_combout ),
	.readdata_17(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[17]~q ),
	.src_data_121(\mm_interconnect_0|rsp_mux|src_data[12]~92_combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux|src_data[11]~96_combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~101_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~107_combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~113_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_009|src_payload~2_combout ),
	.readdata_271(\port_gpio_0|readdata[27]~q ),
	.out_data_buffer_271(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[27]~q ),
	.readdata_281(\port_gpio_0|readdata[28]~q ),
	.out_data_buffer_281(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[28]~q ),
	.readdata_291(\port_gpio_0|readdata[29]~q ),
	.out_data_buffer_291(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[29]~q ),
	.readdata_301(\port_gpio_0|readdata[30]~q ),
	.out_data_buffer_301(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[30]~q ),
	.readdata_31(\port_gpio_0|readdata[31]~q ),
	.out_data_buffer_311(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[31]~q ),
	.readdata_311(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|readdata[31]~q ),
	.debug_reset_request(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_oci_debug|resetrequest~q ),
	.src_payload13(\mm_interconnect_0|cmd_mux_009|src_payload~3_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_009|src_payload~4_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_009|src_payload~5_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_009|src_payload~6_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_009|src_data[33]~combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_009|src_payload~7_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_009|src_payload~8_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_009|src_data[34]~combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_009|src_payload~9_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_009|src_payload~10_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_009|src_payload~11_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_009|src_payload~12_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_009|src_payload~13_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_009|src_payload~14_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_009|src_payload~15_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_009|src_payload~16_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_009|src_payload~17_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_009|src_payload~18_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_009|src_payload~19_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_009|src_data[35]~combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_009|src_payload~20_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_009|src_payload~21_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_009|src_payload~22_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_009|src_payload~23_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_009|src_payload~24_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_009|src_payload~25_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_009|src_payload~26_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_009|src_payload~27_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_009|src_payload~28_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_009|src_payload~29_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_009|src_payload~30_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_009|src_payload~31_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_009|src_payload~32_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ));

niosII_niosII_adc_0 adc_0(
	.wire_pll7_clk_0(\sys_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_4(\cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.sclk(\adc_0|ADC_CTRL|sclk~q ),
	.cs_n(\adc_0|ADC_CTRL|cs_n~2_combout ),
	.addr_shift_reg_5(\adc_0|ADC_CTRL|addr_shift_reg[5]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.mem_used_1(\mm_interconnect_0|adc_0_adc_slave_agent_rsp_fifo|mem_used[1]~q ),
	.Equal3(\mm_interconnect_0|router|Equal3~6_combout ),
	.m0_read(\mm_interconnect_0|adc_0_adc_slave_agent|m0_read~combout ),
	.m0_write(\mm_interconnect_0|timer_0_s1_agent|m0_write~0_combout ),
	.read_mux_out(\timer_0|read_mux_out~0_combout ),
	.d_writedata_0(\cpu|cpu|d_writedata[0]~q ),
	.always0(\adc_0|always0~1_combout ),
	.waitrequest(\adc_0|waitrequest~0_combout ),
	.Equal6(\timer_0|Equal6~1_combout ),
	.av_readdata_pre_0(\mm_interconnect_0|adc_0_adc_slave_translator|av_readdata_pre[0]~0_combout ),
	.readdata_0(\adc_0|readdata[0]~4_combout ),
	.readdata_1(\adc_0|readdata[1]~9_combout ),
	.readdata_2(\adc_0|readdata[2]~14_combout ),
	.readdata_3(\adc_0|readdata[3]~19_combout ),
	.readdata_4(\adc_0|readdata[4]~24_combout ),
	.readdata_5(\adc_0|readdata[5]~29_combout ),
	.readdata_6(\adc_0|readdata[6]~34_combout ),
	.readdata_7(\adc_0|readdata[7]~39_combout ),
	.readdata_15(\adc_0|readdata[15]~40_combout ),
	.readdata_11(\adc_0|readdata[11]~45_combout ),
	.readdata_10(\adc_0|readdata[10]~50_combout ),
	.readdata_9(\adc_0|readdata[9]~55_combout ),
	.readdata_8(\adc_0|readdata[8]~60_combout ),
	.write(\mm_interconnect_0|port_sw_avalon_parallel_port_slave_agent_rsp_fifo|write~3_combout ),
	.GND_port(\~GND~combout ),
	.adc_0_dout(\adc_0_dout~input_o ));

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8 .sum_lutc_input = "datac";

assign \port_gpio_0_export[0]~input_o  = port_gpio_0_export[0];

assign \port_gpio_0_export[1]~input_o  = port_gpio_0_export[1];

assign \port_gpio_0_export[2]~input_o  = port_gpio_0_export[2];

assign \port_gpio_0_export[3]~input_o  = port_gpio_0_export[3];

assign \port_gpio_0_export[4]~input_o  = port_gpio_0_export[4];

assign \port_gpio_0_export[5]~input_o  = port_gpio_0_export[5];

assign \port_gpio_0_export[6]~input_o  = port_gpio_0_export[6];

assign \port_gpio_0_export[7]~input_o  = port_gpio_0_export[7];

assign \port_gpio_0_export[8]~input_o  = port_gpio_0_export[8];

assign \port_gpio_0_export[9]~input_o  = port_gpio_0_export[9];

assign \port_gpio_0_export[10]~input_o  = port_gpio_0_export[10];

assign \port_gpio_0_export[11]~input_o  = port_gpio_0_export[11];

assign \port_gpio_0_export[12]~input_o  = port_gpio_0_export[12];

assign \port_gpio_0_export[13]~input_o  = port_gpio_0_export[13];

assign \port_gpio_0_export[14]~input_o  = port_gpio_0_export[14];

assign \port_gpio_0_export[15]~input_o  = port_gpio_0_export[15];

assign \port_gpio_0_export[16]~input_o  = port_gpio_0_export[16];

assign \port_gpio_0_export[17]~input_o  = port_gpio_0_export[17];

assign \port_gpio_0_export[18]~input_o  = port_gpio_0_export[18];

assign \port_gpio_0_export[19]~input_o  = port_gpio_0_export[19];

assign \port_gpio_0_export[20]~input_o  = port_gpio_0_export[20];

assign \port_gpio_0_export[21]~input_o  = port_gpio_0_export[21];

assign \port_gpio_0_export[22]~input_o  = port_gpio_0_export[22];

assign \port_gpio_0_export[23]~input_o  = port_gpio_0_export[23];

assign \port_gpio_0_export[24]~input_o  = port_gpio_0_export[24];

assign \port_gpio_0_export[25]~input_o  = port_gpio_0_export[25];

assign \port_gpio_0_export[26]~input_o  = port_gpio_0_export[26];

assign \port_gpio_0_export[27]~input_o  = port_gpio_0_export[27];

assign \port_gpio_0_export[28]~input_o  = port_gpio_0_export[28];

assign \port_gpio_0_export[29]~input_o  = port_gpio_0_export[29];

assign \port_gpio_0_export[30]~input_o  = port_gpio_0_export[30];

assign \port_gpio_0_export[31]~input_o  = port_gpio_0_export[31];

assign \sdram_dq[0]~input_o  = sdram_dq[0];

assign \sdram_dq[1]~input_o  = sdram_dq[1];

assign \sdram_dq[2]~input_o  = sdram_dq[2];

assign \sdram_dq[3]~input_o  = sdram_dq[3];

assign \sdram_dq[4]~input_o  = sdram_dq[4];

assign \sdram_dq[5]~input_o  = sdram_dq[5];

assign \sdram_dq[6]~input_o  = sdram_dq[6];

assign \sdram_dq[7]~input_o  = sdram_dq[7];

assign \sdram_dq[8]~input_o  = sdram_dq[8];

assign \sdram_dq[9]~input_o  = sdram_dq[9];

assign \sdram_dq[10]~input_o  = sdram_dq[10];

assign \sdram_dq[11]~input_o  = sdram_dq[11];

assign \sdram_dq[12]~input_o  = sdram_dq[12];

assign \sdram_dq[13]~input_o  = sdram_dq[13];

assign \sdram_dq[14]~input_o  = sdram_dq[14];

assign \sdram_dq[15]~input_o  = sdram_dq[15];

assign \clk_clk~input_o  = clk_clk;

assign \reset_reset_n~input_o  = reset_reset_n;

assign \port_sw_export[0]~input_o  = port_sw_export[0];

assign \port_key_export[0]~input_o  = port_key_export[0];

assign \port_sw_export[1]~input_o  = port_sw_export[1];

assign \port_key_export[1]~input_o  = port_key_export[1];

assign \port_sw_export[2]~input_o  = port_sw_export[2];

assign \port_sw_export[3]~input_o  = port_sw_export[3];

assign \adc_0_dout~input_o  = adc_0_dout;

assign \epcs_data0~input_o  = epcs_data0;

assign \rs232_0_RXD~input_o  = rs232_0_RXD;

assign \rs232_1_RXD~input_o  = rs232_1_RXD;

assign adc_0_sclk = ~ \adc_0|ADC_CTRL|sclk~q ;

assign adc_0_cs_n = ~ \adc_0|ADC_CTRL|cs_n~2_combout ;

assign adc_0_din = \adc_0|ADC_CTRL|addr_shift_reg[5]~q ;

assign epcs_dclk = \epcs|the_niosII_epcs_sub|SCLK_reg~q ;

assign epcs_sce = \epcs|the_niosII_epcs_sub|SS_n~0_combout ;

assign epcs_sdo = \epcs|the_niosII_epcs_sub|shift_reg[7]~q ;

assign port_led_export[0] = \port_led|data_out[0]~q ;

assign port_led_export[1] = \port_led|data_out[1]~q ;

assign port_led_export[2] = \port_led|data_out[2]~q ;

assign port_led_export[3] = \port_led|data_out[3]~q ;

assign port_led_export[4] = \port_led|data_out[4]~q ;

assign port_led_export[5] = \port_led|data_out[5]~q ;

assign port_led_export[6] = \port_led|data_out[6]~q ;

assign port_led_export[7] = \port_led|data_out[7]~q ;

assign ram_clk_clk = \sys_pll|sd1|wire_pll7_clk[1] ;

assign rs232_0_TXD = \rs232_0|RS232_Out_Serializer|serial_data_out~q ;

assign rs232_1_TXD = \rs232_1|RS232_Out_Serializer|serial_data_out~q ;

assign sdram_addr[0] = \sdram|m_addr[0]~q ;

assign sdram_addr[1] = \sdram|m_addr[1]~q ;

assign sdram_addr[2] = \sdram|m_addr[2]~q ;

assign sdram_addr[3] = \sdram|m_addr[3]~q ;

assign sdram_addr[4] = \sdram|m_addr[4]~q ;

assign sdram_addr[5] = \sdram|m_addr[5]~q ;

assign sdram_addr[6] = \sdram|m_addr[6]~q ;

assign sdram_addr[7] = \sdram|m_addr[7]~q ;

assign sdram_addr[8] = \sdram|m_addr[8]~q ;

assign sdram_addr[9] = \sdram|m_addr[9]~q ;

assign sdram_addr[10] = \sdram|m_addr[10]~q ;

assign sdram_addr[11] = \sdram|m_addr[11]~q ;

assign sdram_addr[12] = \sdram|m_addr[12]~q ;

assign sdram_ba[0] = \sdram|m_bank[0]~q ;

assign sdram_ba[1] = \sdram|m_bank[1]~q ;

assign sdram_cas_n = ~ \sdram|m_cmd[1]~q ;

assign sdram_cke = vcc;

assign sdram_cs_n = ~ \sdram|m_cmd[3]~q ;

assign sdram_dqm[0] = \sdram|m_dqm[0]~q ;

assign sdram_dqm[1] = \sdram|m_dqm[1]~q ;

assign sdram_ras_n = ~ \sdram|m_cmd[2]~q ;

assign sdram_we_n = ~ \sdram|m_cmd[0]~q ;

cycloneive_io_obuf \port_gpio_0_export[0]~output (
	.i(\port_gpio_0|data_out[0]~q ),
	.oe(\port_gpio_0|direction[0]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[0]),
	.obar());
defparam \port_gpio_0_export[0]~output .bus_hold = "false";
defparam \port_gpio_0_export[0]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[1]~output (
	.i(\port_gpio_0|data_out[1]~q ),
	.oe(\port_gpio_0|direction[1]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[1]),
	.obar());
defparam \port_gpio_0_export[1]~output .bus_hold = "false";
defparam \port_gpio_0_export[1]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[2]~output (
	.i(\port_gpio_0|data_out[2]~q ),
	.oe(\port_gpio_0|direction[2]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[2]),
	.obar());
defparam \port_gpio_0_export[2]~output .bus_hold = "false";
defparam \port_gpio_0_export[2]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[3]~output (
	.i(\port_gpio_0|data_out[3]~q ),
	.oe(\port_gpio_0|direction[3]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[3]),
	.obar());
defparam \port_gpio_0_export[3]~output .bus_hold = "false";
defparam \port_gpio_0_export[3]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[4]~output (
	.i(\port_gpio_0|data_out[4]~q ),
	.oe(\port_gpio_0|direction[4]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[4]),
	.obar());
defparam \port_gpio_0_export[4]~output .bus_hold = "false";
defparam \port_gpio_0_export[4]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[5]~output (
	.i(\port_gpio_0|data_out[5]~q ),
	.oe(\port_gpio_0|direction[5]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[5]),
	.obar());
defparam \port_gpio_0_export[5]~output .bus_hold = "false";
defparam \port_gpio_0_export[5]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[6]~output (
	.i(\port_gpio_0|data_out[6]~q ),
	.oe(\port_gpio_0|direction[6]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[6]),
	.obar());
defparam \port_gpio_0_export[6]~output .bus_hold = "false";
defparam \port_gpio_0_export[6]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[7]~output (
	.i(\port_gpio_0|data_out[7]~q ),
	.oe(\port_gpio_0|direction[7]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[7]),
	.obar());
defparam \port_gpio_0_export[7]~output .bus_hold = "false";
defparam \port_gpio_0_export[7]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[8]~output (
	.i(\port_gpio_0|data_out[8]~q ),
	.oe(\port_gpio_0|direction[8]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[8]),
	.obar());
defparam \port_gpio_0_export[8]~output .bus_hold = "false";
defparam \port_gpio_0_export[8]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[9]~output (
	.i(\port_gpio_0|data_out[9]~q ),
	.oe(\port_gpio_0|direction[9]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[9]),
	.obar());
defparam \port_gpio_0_export[9]~output .bus_hold = "false";
defparam \port_gpio_0_export[9]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[10]~output (
	.i(\port_gpio_0|data_out[10]~q ),
	.oe(\port_gpio_0|direction[10]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[10]),
	.obar());
defparam \port_gpio_0_export[10]~output .bus_hold = "false";
defparam \port_gpio_0_export[10]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[11]~output (
	.i(\port_gpio_0|data_out[11]~q ),
	.oe(\port_gpio_0|direction[11]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[11]),
	.obar());
defparam \port_gpio_0_export[11]~output .bus_hold = "false";
defparam \port_gpio_0_export[11]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[12]~output (
	.i(\port_gpio_0|data_out[12]~q ),
	.oe(\port_gpio_0|direction[12]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[12]),
	.obar());
defparam \port_gpio_0_export[12]~output .bus_hold = "false";
defparam \port_gpio_0_export[12]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[13]~output (
	.i(\port_gpio_0|data_out[13]~q ),
	.oe(\port_gpio_0|direction[13]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[13]),
	.obar());
defparam \port_gpio_0_export[13]~output .bus_hold = "false";
defparam \port_gpio_0_export[13]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[14]~output (
	.i(\port_gpio_0|data_out[14]~q ),
	.oe(\port_gpio_0|direction[14]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[14]),
	.obar());
defparam \port_gpio_0_export[14]~output .bus_hold = "false";
defparam \port_gpio_0_export[14]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[15]~output (
	.i(\port_gpio_0|data_out[15]~q ),
	.oe(\port_gpio_0|direction[15]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[15]),
	.obar());
defparam \port_gpio_0_export[15]~output .bus_hold = "false";
defparam \port_gpio_0_export[15]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[16]~output (
	.i(\port_gpio_0|data_out[16]~q ),
	.oe(\port_gpio_0|direction[16]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[16]),
	.obar());
defparam \port_gpio_0_export[16]~output .bus_hold = "false";
defparam \port_gpio_0_export[16]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[17]~output (
	.i(\port_gpio_0|data_out[17]~q ),
	.oe(\port_gpio_0|direction[17]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[17]),
	.obar());
defparam \port_gpio_0_export[17]~output .bus_hold = "false";
defparam \port_gpio_0_export[17]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[18]~output (
	.i(\port_gpio_0|data_out[18]~q ),
	.oe(\port_gpio_0|direction[18]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[18]),
	.obar());
defparam \port_gpio_0_export[18]~output .bus_hold = "false";
defparam \port_gpio_0_export[18]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[19]~output (
	.i(\port_gpio_0|data_out[19]~q ),
	.oe(\port_gpio_0|direction[19]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[19]),
	.obar());
defparam \port_gpio_0_export[19]~output .bus_hold = "false";
defparam \port_gpio_0_export[19]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[20]~output (
	.i(\port_gpio_0|data_out[20]~q ),
	.oe(\port_gpio_0|direction[20]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[20]),
	.obar());
defparam \port_gpio_0_export[20]~output .bus_hold = "false";
defparam \port_gpio_0_export[20]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[21]~output (
	.i(\port_gpio_0|data_out[21]~q ),
	.oe(\port_gpio_0|direction[21]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[21]),
	.obar());
defparam \port_gpio_0_export[21]~output .bus_hold = "false";
defparam \port_gpio_0_export[21]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[22]~output (
	.i(\port_gpio_0|data_out[22]~q ),
	.oe(\port_gpio_0|direction[22]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[22]),
	.obar());
defparam \port_gpio_0_export[22]~output .bus_hold = "false";
defparam \port_gpio_0_export[22]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[23]~output (
	.i(\port_gpio_0|data_out[23]~q ),
	.oe(\port_gpio_0|direction[23]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[23]),
	.obar());
defparam \port_gpio_0_export[23]~output .bus_hold = "false";
defparam \port_gpio_0_export[23]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[24]~output (
	.i(\port_gpio_0|data_out[24]~q ),
	.oe(\port_gpio_0|direction[24]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[24]),
	.obar());
defparam \port_gpio_0_export[24]~output .bus_hold = "false";
defparam \port_gpio_0_export[24]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[25]~output (
	.i(\port_gpio_0|data_out[25]~q ),
	.oe(\port_gpio_0|direction[25]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[25]),
	.obar());
defparam \port_gpio_0_export[25]~output .bus_hold = "false";
defparam \port_gpio_0_export[25]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[26]~output (
	.i(\port_gpio_0|data_out[26]~q ),
	.oe(\port_gpio_0|direction[26]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[26]),
	.obar());
defparam \port_gpio_0_export[26]~output .bus_hold = "false";
defparam \port_gpio_0_export[26]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[27]~output (
	.i(\port_gpio_0|data_out[27]~q ),
	.oe(\port_gpio_0|direction[27]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[27]),
	.obar());
defparam \port_gpio_0_export[27]~output .bus_hold = "false";
defparam \port_gpio_0_export[27]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[28]~output (
	.i(\port_gpio_0|data_out[28]~q ),
	.oe(\port_gpio_0|direction[28]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[28]),
	.obar());
defparam \port_gpio_0_export[28]~output .bus_hold = "false";
defparam \port_gpio_0_export[28]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[29]~output (
	.i(\port_gpio_0|data_out[29]~q ),
	.oe(\port_gpio_0|direction[29]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[29]),
	.obar());
defparam \port_gpio_0_export[29]~output .bus_hold = "false";
defparam \port_gpio_0_export[29]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[30]~output (
	.i(\port_gpio_0|data_out[30]~q ),
	.oe(\port_gpio_0|direction[30]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[30]),
	.obar());
defparam \port_gpio_0_export[30]~output .bus_hold = "false";
defparam \port_gpio_0_export[30]~output .open_drain_output = "false";

cycloneive_io_obuf \port_gpio_0_export[31]~output (
	.i(\port_gpio_0|data_out[31]~q ),
	.oe(\port_gpio_0|direction[31]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(port_gpio_0_export[31]),
	.obar());
defparam \port_gpio_0_export[31]~output .bus_hold = "false";
defparam \port_gpio_0_export[31]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[0]~output (
	.i(\sdram|m_data[0]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[0]),
	.obar());
defparam \sdram_dq[0]~output .bus_hold = "false";
defparam \sdram_dq[0]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[1]~output (
	.i(\sdram|m_data[1]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[1]),
	.obar());
defparam \sdram_dq[1]~output .bus_hold = "false";
defparam \sdram_dq[1]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[2]~output (
	.i(\sdram|m_data[2]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[2]),
	.obar());
defparam \sdram_dq[2]~output .bus_hold = "false";
defparam \sdram_dq[2]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[3]~output (
	.i(\sdram|m_data[3]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[3]),
	.obar());
defparam \sdram_dq[3]~output .bus_hold = "false";
defparam \sdram_dq[3]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[4]~output (
	.i(\sdram|m_data[4]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[4]),
	.obar());
defparam \sdram_dq[4]~output .bus_hold = "false";
defparam \sdram_dq[4]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[5]~output (
	.i(\sdram|m_data[5]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[5]),
	.obar());
defparam \sdram_dq[5]~output .bus_hold = "false";
defparam \sdram_dq[5]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[6]~output (
	.i(\sdram|m_data[6]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[6]),
	.obar());
defparam \sdram_dq[6]~output .bus_hold = "false";
defparam \sdram_dq[6]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[7]~output (
	.i(\sdram|m_data[7]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[7]),
	.obar());
defparam \sdram_dq[7]~output .bus_hold = "false";
defparam \sdram_dq[7]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[8]~output (
	.i(\sdram|m_data[8]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[8]),
	.obar());
defparam \sdram_dq[8]~output .bus_hold = "false";
defparam \sdram_dq[8]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[9]~output (
	.i(\sdram|m_data[9]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[9]),
	.obar());
defparam \sdram_dq[9]~output .bus_hold = "false";
defparam \sdram_dq[9]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[10]~output (
	.i(\sdram|m_data[10]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[10]),
	.obar());
defparam \sdram_dq[10]~output .bus_hold = "false";
defparam \sdram_dq[10]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[11]~output (
	.i(\sdram|m_data[11]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[11]),
	.obar());
defparam \sdram_dq[11]~output .bus_hold = "false";
defparam \sdram_dq[11]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[12]~output (
	.i(\sdram|m_data[12]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[12]),
	.obar());
defparam \sdram_dq[12]~output .bus_hold = "false";
defparam \sdram_dq[12]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[13]~output (
	.i(\sdram|m_data[13]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[13]),
	.obar());
defparam \sdram_dq[13]~output .bus_hold = "false";
defparam \sdram_dq[13]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[14]~output (
	.i(\sdram|m_data[14]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[14]),
	.obar());
defparam \sdram_dq[14]~output .bus_hold = "false";
defparam \sdram_dq[14]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_dq[15]~output (
	.i(\sdram|m_data[15]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_dq[15]),
	.obar());
defparam \sdram_dq[15]~output .bus_hold = "false";
defparam \sdram_dq[15]~output .open_drain_output = "false";

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\~GND~combout ),
	.datad(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7_combout ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 (
	.dataa(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|ir_out[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10 .lut_mask = 16'hFFB8;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8 .lut_mask = 16'hF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .lut_mask = 16'h8B8B;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 (
	.dataa(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|ir_out[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\jtag|niosII_jtag_alt_jtag_atlantic|tdo~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~7_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~8 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~7 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~8 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~11 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~13 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~13 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~15_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~16 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~15 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~15 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~16 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~17 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~17 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~19_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 16'hFBFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 16'h27FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~6 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 16'hC5C5;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 16'hD77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 16'hDEDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .lut_mask = 16'hD77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .lut_mask = 16'hFFFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23 .lut_mask = 16'hFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 .lut_mask = 16'hFF6F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .lut_mask = 16'hFFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .lut_mask = 16'hBF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 16'hFFBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 16'hFFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(\jtag|niosII_jtag_alt_jtag_atlantic|tdo~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datab(\cpu|cpu|the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";

endmodule

module niosII_altera_irq_clock_crosser (
	wire_pll7_clk_0,
	r_sync_rst,
	dreg_1,
	av_irq)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
output 	dreg_1;
input 	av_irq;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_std_synchronizer_bundle_1 sync(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.dreg_1(dreg_1),
	.av_irq(av_irq));

endmodule

module niosII_altera_irq_clock_crosser_1 (
	wire_pll7_clk_0,
	r_sync_rst,
	dreg_1,
	irq_reg)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
output 	dreg_1;
input 	irq_reg;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_std_synchronizer_bundle sync(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.dreg_1(dreg_1),
	.irq_reg(irq_reg));

endmodule

module niosII_altera_std_synchronizer_bundle (
	wire_pll7_clk_0,
	r_sync_rst,
	dreg_1,
	irq_reg)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
output 	dreg_1;
input 	irq_reg;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_std_synchronizer \sync[0].u (
	.clk(wire_pll7_clk_0),
	.reset_n(r_sync_rst),
	.dreg_1(dreg_1),
	.din(irq_reg));

endmodule

module niosII_altera_std_synchronizer (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_bundle_1 (
	wire_pll7_clk_0,
	r_sync_rst,
	dreg_1,
	av_irq)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
output 	dreg_1;
input 	av_irq;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_std_synchronizer_1 \sync[0].u (
	.clk(wire_pll7_clk_0),
	.reset_n(r_sync_rst),
	.dreg_1(dreg_1),
	.din(av_irq));

endmodule

module niosII_altera_std_synchronizer_1 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module niosII_altera_reset_controller (
	wire_pll7_clk_0,
	r_sync_rst1,
	r_early_rst1,
	altera_reset_synchronizer_int_chain_1,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	r_sync_rst1;
output 	r_early_rst1;
output 	altera_reset_synchronizer_int_chain_1;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


niosII_altera_reset_synchronizer_5 alt_rst_sync_uq1(
	.clk(wire_pll7_clk_0),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.reset_reset_n(reset_reset_n));

niosII_altera_reset_synchronizer_4 alt_rst_req_sync_uq1(
	.clk(wire_pll7_clk_0),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1));

dffeas r_sync_rst(
	.clk(wire_pll7_clk_0),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(wire_pll7_clk_0),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(wire_pll7_clk_0),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.cout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 16'h5555;
defparam \altera_reset_synchronizer_int_chain[4]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[3]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.cout());
defparam \r_sync_rst_chain~1 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~1 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[2] (
	.clk(wire_pll7_clk_0),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.cout());
defparam \r_sync_rst_chain~0 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~0 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[1] (
	.clk(wire_pll7_clk_0),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(\altera_reset_synchronizer_int_chain[4]~q ),
	.datab(r_sync_rst1),
	.datac(gnd),
	.datad(\r_sync_rst_chain[1]~q ),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEEFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hAAFF;
defparam \always2~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_reset_controller_1 (
	wire_pll7_clk_0,
	r_sync_rst1,
	resetrequest,
	r_early_rst1,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	r_sync_rst1;
input 	resetrequest;
output 	r_early_rst1;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \merged_reset~0_combout ;
wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


niosII_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.clk(wire_pll7_clk_0),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ));

niosII_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.clk(wire_pll7_clk_0),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.merged_reset(\merged_reset~0_combout ));

cycloneive_lcell_comb \merged_reset~0 (
	.dataa(resetrequest),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_reset_n),
	.cin(gnd),
	.combout(\merged_reset~0_combout ),
	.cout());
defparam \merged_reset~0 .lut_mask = 16'hAAFF;
defparam \merged_reset~0 .sum_lutc_input = "datac";

dffeas r_sync_rst(
	.clk(wire_pll7_clk_0),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(wire_pll7_clk_0),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(wire_pll7_clk_0),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.cout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 16'h5555;
defparam \altera_reset_synchronizer_int_chain[4]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(wire_pll7_clk_0),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[3]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.cout());
defparam \r_sync_rst_chain~1 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~1 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[2] (
	.clk(wire_pll7_clk_0),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.cout());
defparam \r_sync_rst_chain~0 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~0 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[1] (
	.clk(wire_pll7_clk_0),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(\altera_reset_synchronizer_int_chain[4]~q ),
	.datab(r_sync_rst1),
	.datac(gnd),
	.datad(\r_sync_rst_chain[1]~q ),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEEFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hAAFF;
defparam \always2~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_reset_synchronizer (
	clk,
	altera_reset_synchronizer_int_chain_out1)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.cout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 16'h0000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module niosII_altera_reset_synchronizer_1 (
	clk,
	altera_reset_synchronizer_int_chain_out1,
	merged_reset)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;
input 	merged_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module niosII_altera_reset_controller_2 (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module niosII_altera_reset_synchronizer_3 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module niosII_altera_reset_synchronizer_4 (
	clk,
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.cout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 16'h0000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module niosII_altera_reset_synchronizer_5 (
	clk,
	altera_reset_synchronizer_int_chain_out1,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module niosII_niosII_adc_0 (
	wire_pll7_clk_0,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	sclk,
	cs_n,
	addr_shift_reg_5,
	r_sync_rst,
	mem_used_1,
	Equal3,
	m0_read,
	m0_write,
	read_mux_out,
	d_writedata_0,
	always0,
	waitrequest,
	Equal6,
	av_readdata_pre_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_15,
	readdata_11,
	readdata_10,
	readdata_9,
	readdata_8,
	write,
	GND_port,
	adc_0_dout)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
output 	sclk;
output 	cs_n;
output 	addr_shift_reg_5;
input 	r_sync_rst;
input 	mem_used_1;
input 	Equal3;
input 	m0_read;
input 	m0_write;
input 	read_mux_out;
input 	d_writedata_0;
output 	always0;
output 	waitrequest;
input 	Equal6;
input 	av_readdata_pre_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_15;
output 	readdata_11;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
input 	write;
input 	GND_port;
input 	adc_0_dout;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ADC_CTRL|currState.doneState~q ;
wire \ADC_CTRL|reading6[0]~q ;
wire \ADC_CTRL|reading5[0]~q ;
wire \ADC_CTRL|reading4[0]~q ;
wire \ADC_CTRL|reading7[0]~q ;
wire \ADC_CTRL|reading2[0]~q ;
wire \ADC_CTRL|reading1[0]~q ;
wire \ADC_CTRL|reading0[0]~q ;
wire \ADC_CTRL|reading3[0]~q ;
wire \ADC_CTRL|reading6[1]~q ;
wire \ADC_CTRL|reading5[1]~q ;
wire \ADC_CTRL|reading4[1]~q ;
wire \ADC_CTRL|reading7[1]~q ;
wire \ADC_CTRL|reading2[1]~q ;
wire \ADC_CTRL|reading1[1]~q ;
wire \ADC_CTRL|reading0[1]~q ;
wire \ADC_CTRL|reading3[1]~q ;
wire \ADC_CTRL|reading6[2]~q ;
wire \ADC_CTRL|reading5[2]~q ;
wire \ADC_CTRL|reading4[2]~q ;
wire \ADC_CTRL|reading7[2]~q ;
wire \ADC_CTRL|reading2[2]~q ;
wire \ADC_CTRL|reading1[2]~q ;
wire \ADC_CTRL|reading0[2]~q ;
wire \ADC_CTRL|reading3[2]~q ;
wire \ADC_CTRL|reading6[3]~q ;
wire \ADC_CTRL|reading5[3]~q ;
wire \ADC_CTRL|reading4[3]~q ;
wire \ADC_CTRL|reading7[3]~q ;
wire \ADC_CTRL|reading2[3]~q ;
wire \ADC_CTRL|reading1[3]~q ;
wire \ADC_CTRL|reading0[3]~q ;
wire \ADC_CTRL|reading3[3]~q ;
wire \ADC_CTRL|reading6[4]~q ;
wire \ADC_CTRL|reading5[4]~q ;
wire \ADC_CTRL|reading4[4]~q ;
wire \ADC_CTRL|reading7[4]~q ;
wire \ADC_CTRL|reading2[4]~q ;
wire \ADC_CTRL|reading1[4]~q ;
wire \ADC_CTRL|reading0[4]~q ;
wire \ADC_CTRL|reading3[4]~q ;
wire \ADC_CTRL|reading6[5]~q ;
wire \ADC_CTRL|reading5[5]~q ;
wire \ADC_CTRL|reading4[5]~q ;
wire \ADC_CTRL|reading7[5]~q ;
wire \ADC_CTRL|reading2[5]~q ;
wire \ADC_CTRL|reading1[5]~q ;
wire \ADC_CTRL|reading0[5]~q ;
wire \ADC_CTRL|reading3[5]~q ;
wire \ADC_CTRL|reading6[6]~q ;
wire \ADC_CTRL|reading5[6]~q ;
wire \ADC_CTRL|reading4[6]~q ;
wire \ADC_CTRL|reading7[6]~q ;
wire \ADC_CTRL|reading2[6]~q ;
wire \ADC_CTRL|reading1[6]~q ;
wire \ADC_CTRL|reading0[6]~q ;
wire \ADC_CTRL|reading3[6]~q ;
wire \ADC_CTRL|reading6[7]~q ;
wire \ADC_CTRL|reading5[7]~q ;
wire \ADC_CTRL|reading4[7]~q ;
wire \ADC_CTRL|reading7[7]~q ;
wire \ADC_CTRL|reading2[7]~q ;
wire \ADC_CTRL|reading1[7]~q ;
wire \ADC_CTRL|reading0[7]~q ;
wire \ADC_CTRL|reading3[7]~q ;
wire \ADC_CTRL|reading6[11]~q ;
wire \ADC_CTRL|reading5[11]~q ;
wire \ADC_CTRL|reading4[11]~q ;
wire \ADC_CTRL|reading7[11]~q ;
wire \ADC_CTRL|reading2[11]~q ;
wire \ADC_CTRL|reading1[11]~q ;
wire \ADC_CTRL|reading0[11]~q ;
wire \ADC_CTRL|reading3[11]~q ;
wire \ADC_CTRL|reading6[10]~q ;
wire \ADC_CTRL|reading5[10]~q ;
wire \ADC_CTRL|reading4[10]~q ;
wire \ADC_CTRL|reading7[10]~q ;
wire \ADC_CTRL|reading2[10]~q ;
wire \ADC_CTRL|reading1[10]~q ;
wire \ADC_CTRL|reading0[10]~q ;
wire \ADC_CTRL|reading3[10]~q ;
wire \ADC_CTRL|reading6[9]~q ;
wire \ADC_CTRL|reading5[9]~q ;
wire \ADC_CTRL|reading4[9]~q ;
wire \ADC_CTRL|reading7[9]~q ;
wire \ADC_CTRL|reading2[9]~q ;
wire \ADC_CTRL|reading1[9]~q ;
wire \ADC_CTRL|reading0[9]~q ;
wire \ADC_CTRL|reading3[9]~q ;
wire \ADC_CTRL|reading6[8]~q ;
wire \ADC_CTRL|reading5[8]~q ;
wire \ADC_CTRL|reading4[8]~q ;
wire \ADC_CTRL|reading7[8]~q ;
wire \ADC_CTRL|reading2[8]~q ;
wire \ADC_CTRL|reading1[8]~q ;
wire \ADC_CTRL|reading0[8]~q ;
wire \ADC_CTRL|reading3[8]~q ;
wire \always0~0_combout ;
wire \auto_run~0_combout ;
wire \auto_run~q ;
wire \go~0_combout ;
wire \go~1_combout ;
wire \go~q ;
wire \values[6][0]~q ;
wire \values[5][0]~q ;
wire \values[4][0]~q ;
wire \readdata[0]~0_combout ;
wire \values[7][0]~q ;
wire \readdata[0]~1_combout ;
wire \values[2][0]~q ;
wire \values[1][0]~q ;
wire \values[0][0]~q ;
wire \readdata[0]~2_combout ;
wire \values[3][0]~q ;
wire \readdata[0]~3_combout ;
wire \values[6][1]~q ;
wire \values[5][1]~q ;
wire \values[4][1]~q ;
wire \readdata[1]~5_combout ;
wire \values[7][1]~q ;
wire \readdata[1]~6_combout ;
wire \values[2][1]~q ;
wire \values[1][1]~q ;
wire \values[0][1]~q ;
wire \readdata[1]~7_combout ;
wire \values[3][1]~q ;
wire \readdata[1]~8_combout ;
wire \values[6][2]~q ;
wire \values[5][2]~q ;
wire \values[4][2]~q ;
wire \readdata[2]~10_combout ;
wire \values[7][2]~q ;
wire \readdata[2]~11_combout ;
wire \values[2][2]~q ;
wire \values[1][2]~q ;
wire \values[0][2]~q ;
wire \readdata[2]~12_combout ;
wire \values[3][2]~q ;
wire \readdata[2]~13_combout ;
wire \values[6][3]~q ;
wire \values[5][3]~q ;
wire \values[4][3]~q ;
wire \readdata[3]~15_combout ;
wire \values[7][3]~q ;
wire \readdata[3]~16_combout ;
wire \values[2][3]~q ;
wire \values[1][3]~q ;
wire \values[0][3]~q ;
wire \readdata[3]~17_combout ;
wire \values[3][3]~q ;
wire \readdata[3]~18_combout ;
wire \values[6][4]~q ;
wire \values[5][4]~q ;
wire \values[4][4]~q ;
wire \readdata[4]~20_combout ;
wire \values[7][4]~q ;
wire \readdata[4]~21_combout ;
wire \values[2][4]~q ;
wire \values[1][4]~q ;
wire \values[0][4]~q ;
wire \readdata[4]~22_combout ;
wire \values[3][4]~q ;
wire \readdata[4]~23_combout ;
wire \values[6][5]~q ;
wire \values[5][5]~q ;
wire \values[4][5]~q ;
wire \readdata[5]~25_combout ;
wire \values[7][5]~q ;
wire \readdata[5]~26_combout ;
wire \values[2][5]~q ;
wire \values[1][5]~q ;
wire \values[0][5]~q ;
wire \readdata[5]~27_combout ;
wire \values[3][5]~q ;
wire \readdata[5]~28_combout ;
wire \values[6][6]~q ;
wire \values[5][6]~q ;
wire \values[4][6]~q ;
wire \readdata[6]~30_combout ;
wire \values[7][6]~q ;
wire \readdata[6]~31_combout ;
wire \values[2][6]~q ;
wire \values[1][6]~q ;
wire \values[0][6]~q ;
wire \readdata[6]~32_combout ;
wire \values[3][6]~q ;
wire \readdata[6]~33_combout ;
wire \values[6][7]~q ;
wire \values[5][7]~q ;
wire \values[4][7]~q ;
wire \readdata[7]~35_combout ;
wire \values[7][7]~q ;
wire \readdata[7]~36_combout ;
wire \values[2][7]~q ;
wire \values[1][7]~q ;
wire \values[0][7]~q ;
wire \readdata[7]~37_combout ;
wire \values[3][7]~q ;
wire \readdata[7]~38_combout ;
wire \always1~0_combout ;
wire \Decoder0~0_combout ;
wire \refresh~0_combout ;
wire \refresh[5]~q ;
wire \Decoder0~1_combout ;
wire \refresh~1_combout ;
wire \refresh[6]~q ;
wire \Decoder0~2_combout ;
wire \refresh~2_combout ;
wire \refresh[4]~q ;
wire \Mux0~0_combout ;
wire \Decoder0~3_combout ;
wire \refresh~3_combout ;
wire \refresh[7]~q ;
wire \Mux0~1_combout ;
wire \Decoder0~4_combout ;
wire \refresh~4_combout ;
wire \refresh[2]~q ;
wire \Decoder0~5_combout ;
wire \refresh~5_combout ;
wire \refresh[1]~q ;
wire \Decoder0~6_combout ;
wire \refresh~6_combout ;
wire \refresh[0]~q ;
wire \Mux0~2_combout ;
wire \Decoder0~7_combout ;
wire \refresh~7_combout ;
wire \refresh[3]~q ;
wire \Mux0~3_combout ;
wire \values[6][11]~q ;
wire \values[5][11]~q ;
wire \values[4][11]~q ;
wire \readdata[11]~41_combout ;
wire \values[7][11]~q ;
wire \readdata[11]~42_combout ;
wire \values[2][11]~q ;
wire \values[1][11]~q ;
wire \values[0][11]~q ;
wire \readdata[11]~43_combout ;
wire \values[3][11]~q ;
wire \readdata[11]~44_combout ;
wire \values[6][10]~q ;
wire \values[5][10]~q ;
wire \values[4][10]~q ;
wire \readdata[10]~46_combout ;
wire \values[7][10]~q ;
wire \readdata[10]~47_combout ;
wire \values[2][10]~q ;
wire \values[1][10]~q ;
wire \values[0][10]~q ;
wire \readdata[10]~48_combout ;
wire \values[3][10]~q ;
wire \readdata[10]~49_combout ;
wire \values[6][9]~q ;
wire \values[5][9]~q ;
wire \values[4][9]~q ;
wire \readdata[9]~51_combout ;
wire \values[7][9]~q ;
wire \readdata[9]~52_combout ;
wire \values[2][9]~q ;
wire \values[1][9]~q ;
wire \values[0][9]~q ;
wire \readdata[9]~53_combout ;
wire \values[3][9]~q ;
wire \readdata[9]~54_combout ;
wire \values[6][8]~q ;
wire \values[5][8]~q ;
wire \values[4][8]~q ;
wire \readdata[8]~56_combout ;
wire \values[7][8]~q ;
wire \readdata[8]~57_combout ;
wire \values[2][8]~q ;
wire \values[1][8]~q ;
wire \values[0][8]~q ;
wire \readdata[8]~58_combout ;
wire \values[3][8]~q ;
wire \readdata[8]~59_combout ;


niosII_altera_up_avalon_adv_adc ADC_CTRL(
	.clock(wire_pll7_clk_0),
	.go(\go~q ),
	.sclk1(sclk),
	.cs_n(cs_n),
	.addr_shift_reg_5(addr_shift_reg_5),
	.r_sync_rst(r_sync_rst),
	.currStatedoneState(\ADC_CTRL|currState.doneState~q ),
	.reading6_0(\ADC_CTRL|reading6[0]~q ),
	.reading5_0(\ADC_CTRL|reading5[0]~q ),
	.reading4_0(\ADC_CTRL|reading4[0]~q ),
	.reading7_0(\ADC_CTRL|reading7[0]~q ),
	.reading2_0(\ADC_CTRL|reading2[0]~q ),
	.reading1_0(\ADC_CTRL|reading1[0]~q ),
	.reading0_0(\ADC_CTRL|reading0[0]~q ),
	.reading3_0(\ADC_CTRL|reading3[0]~q ),
	.reading6_1(\ADC_CTRL|reading6[1]~q ),
	.reading5_1(\ADC_CTRL|reading5[1]~q ),
	.reading4_1(\ADC_CTRL|reading4[1]~q ),
	.reading7_1(\ADC_CTRL|reading7[1]~q ),
	.reading2_1(\ADC_CTRL|reading2[1]~q ),
	.reading1_1(\ADC_CTRL|reading1[1]~q ),
	.reading0_1(\ADC_CTRL|reading0[1]~q ),
	.reading3_1(\ADC_CTRL|reading3[1]~q ),
	.reading6_2(\ADC_CTRL|reading6[2]~q ),
	.reading5_2(\ADC_CTRL|reading5[2]~q ),
	.reading4_2(\ADC_CTRL|reading4[2]~q ),
	.reading7_2(\ADC_CTRL|reading7[2]~q ),
	.reading2_2(\ADC_CTRL|reading2[2]~q ),
	.reading1_2(\ADC_CTRL|reading1[2]~q ),
	.reading0_2(\ADC_CTRL|reading0[2]~q ),
	.reading3_2(\ADC_CTRL|reading3[2]~q ),
	.reading6_3(\ADC_CTRL|reading6[3]~q ),
	.reading5_3(\ADC_CTRL|reading5[3]~q ),
	.reading4_3(\ADC_CTRL|reading4[3]~q ),
	.reading7_3(\ADC_CTRL|reading7[3]~q ),
	.reading2_3(\ADC_CTRL|reading2[3]~q ),
	.reading1_3(\ADC_CTRL|reading1[3]~q ),
	.reading0_3(\ADC_CTRL|reading0[3]~q ),
	.reading3_3(\ADC_CTRL|reading3[3]~q ),
	.reading6_4(\ADC_CTRL|reading6[4]~q ),
	.reading5_4(\ADC_CTRL|reading5[4]~q ),
	.reading4_4(\ADC_CTRL|reading4[4]~q ),
	.reading7_4(\ADC_CTRL|reading7[4]~q ),
	.reading2_4(\ADC_CTRL|reading2[4]~q ),
	.reading1_4(\ADC_CTRL|reading1[4]~q ),
	.reading0_4(\ADC_CTRL|reading0[4]~q ),
	.reading3_4(\ADC_CTRL|reading3[4]~q ),
	.reading6_5(\ADC_CTRL|reading6[5]~q ),
	.reading5_5(\ADC_CTRL|reading5[5]~q ),
	.reading4_5(\ADC_CTRL|reading4[5]~q ),
	.reading7_5(\ADC_CTRL|reading7[5]~q ),
	.reading2_5(\ADC_CTRL|reading2[5]~q ),
	.reading1_5(\ADC_CTRL|reading1[5]~q ),
	.reading0_5(\ADC_CTRL|reading0[5]~q ),
	.reading3_5(\ADC_CTRL|reading3[5]~q ),
	.reading6_6(\ADC_CTRL|reading6[6]~q ),
	.reading5_6(\ADC_CTRL|reading5[6]~q ),
	.reading4_6(\ADC_CTRL|reading4[6]~q ),
	.reading7_6(\ADC_CTRL|reading7[6]~q ),
	.reading2_6(\ADC_CTRL|reading2[6]~q ),
	.reading1_6(\ADC_CTRL|reading1[6]~q ),
	.reading0_6(\ADC_CTRL|reading0[6]~q ),
	.reading3_6(\ADC_CTRL|reading3[6]~q ),
	.reading6_7(\ADC_CTRL|reading6[7]~q ),
	.reading5_7(\ADC_CTRL|reading5[7]~q ),
	.reading4_7(\ADC_CTRL|reading4[7]~q ),
	.reading7_7(\ADC_CTRL|reading7[7]~q ),
	.reading2_7(\ADC_CTRL|reading2[7]~q ),
	.reading1_7(\ADC_CTRL|reading1[7]~q ),
	.reading0_7(\ADC_CTRL|reading0[7]~q ),
	.reading3_7(\ADC_CTRL|reading3[7]~q ),
	.reading6_11(\ADC_CTRL|reading6[11]~q ),
	.reading5_11(\ADC_CTRL|reading5[11]~q ),
	.reading4_11(\ADC_CTRL|reading4[11]~q ),
	.reading7_11(\ADC_CTRL|reading7[11]~q ),
	.reading2_11(\ADC_CTRL|reading2[11]~q ),
	.reading1_11(\ADC_CTRL|reading1[11]~q ),
	.reading0_11(\ADC_CTRL|reading0[11]~q ),
	.reading3_11(\ADC_CTRL|reading3[11]~q ),
	.reading6_10(\ADC_CTRL|reading6[10]~q ),
	.reading5_10(\ADC_CTRL|reading5[10]~q ),
	.reading4_10(\ADC_CTRL|reading4[10]~q ),
	.reading7_10(\ADC_CTRL|reading7[10]~q ),
	.reading2_10(\ADC_CTRL|reading2[10]~q ),
	.reading1_10(\ADC_CTRL|reading1[10]~q ),
	.reading0_10(\ADC_CTRL|reading0[10]~q ),
	.reading3_10(\ADC_CTRL|reading3[10]~q ),
	.reading6_9(\ADC_CTRL|reading6[9]~q ),
	.reading5_9(\ADC_CTRL|reading5[9]~q ),
	.reading4_9(\ADC_CTRL|reading4[9]~q ),
	.reading7_9(\ADC_CTRL|reading7[9]~q ),
	.reading2_9(\ADC_CTRL|reading2[9]~q ),
	.reading1_9(\ADC_CTRL|reading1[9]~q ),
	.reading0_9(\ADC_CTRL|reading0[9]~q ),
	.reading3_9(\ADC_CTRL|reading3[9]~q ),
	.reading6_8(\ADC_CTRL|reading6[8]~q ),
	.reading5_8(\ADC_CTRL|reading5[8]~q ),
	.reading4_8(\ADC_CTRL|reading4[8]~q ),
	.reading7_8(\ADC_CTRL|reading7[8]~q ),
	.reading2_8(\ADC_CTRL|reading2[8]~q ),
	.reading1_8(\ADC_CTRL|reading1[8]~q ),
	.reading0_8(\ADC_CTRL|reading0[8]~q ),
	.reading3_8(\ADC_CTRL|reading3[8]~q ),
	.dout(adc_0_dout));

cycloneive_lcell_comb \always0~1 (
	.dataa(\go~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_run~q ),
	.cin(gnd),
	.combout(always0),
	.cout());
defparam \always0~1 .lut_mask = 16'hAAFF;
defparam \always0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \waitrequest~0 (
	.dataa(\ADC_CTRL|currState.doneState~q ),
	.datab(\always0~0_combout ),
	.datac(always0),
	.datad(m0_read),
	.cin(gnd),
	.combout(waitrequest),
	.cout());
defparam \waitrequest~0 .lut_mask = 16'hFEFF;
defparam \waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0]~4 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[0]~1_combout ),
	.datac(\readdata[0]~3_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0]~4 .lut_mask = 16'hFAFC;
defparam \readdata[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1]~9 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[1]~6_combout ),
	.datac(\readdata[1]~8_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1]~9 .lut_mask = 16'hFAFC;
defparam \readdata[1]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[2]~14 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[2]~11_combout ),
	.datac(\readdata[2]~13_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2]~14 .lut_mask = 16'hFAFC;
defparam \readdata[2]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3]~19 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[3]~16_combout ),
	.datac(\readdata[3]~18_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3]~19 .lut_mask = 16'hFAFC;
defparam \readdata[3]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[4]~24 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[4]~21_combout ),
	.datac(\readdata[4]~23_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4]~24 .lut_mask = 16'hFAFC;
defparam \readdata[4]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[5]~29 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[5]~26_combout ),
	.datac(\readdata[5]~28_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5]~29 .lut_mask = 16'hFAFC;
defparam \readdata[5]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[6]~34 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[6]~31_combout ),
	.datac(\readdata[6]~33_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6]~34 .lut_mask = 16'hFAFC;
defparam \readdata[6]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[7]~39 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[7]~36_combout ),
	.datac(\readdata[7]~38_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7]~39 .lut_mask = 16'hFAFC;
defparam \readdata[7]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[15]~40 (
	.dataa(\always1~0_combout ),
	.datab(\Mux0~1_combout ),
	.datac(\Mux0~3_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_15),
	.cout());
defparam \readdata[15]~40 .lut_mask = 16'hFAFC;
defparam \readdata[15]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[11]~45 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[11]~42_combout ),
	.datac(\readdata[11]~44_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_11),
	.cout());
defparam \readdata[11]~45 .lut_mask = 16'hFAFC;
defparam \readdata[11]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[10]~50 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[10]~47_combout ),
	.datac(\readdata[10]~49_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_10),
	.cout());
defparam \readdata[10]~50 .lut_mask = 16'hFAFC;
defparam \readdata[10]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[9]~55 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[9]~52_combout ),
	.datac(\readdata[9]~54_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_9),
	.cout());
defparam \readdata[9]~55 .lut_mask = 16'hFAFC;
defparam \readdata[9]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[8]~60 (
	.dataa(av_readdata_pre_0),
	.datab(\readdata[8]~57_combout ),
	.datac(\readdata[8]~59_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(readdata_8),
	.cout());
defparam \readdata[8]~60 .lut_mask = 16'hFAFC;
defparam \readdata[8]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(Equal3),
	.datab(m0_write),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hEEFF;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_run~0 (
	.dataa(d_writedata_0),
	.datab(\auto_run~q ),
	.datac(\always0~0_combout ),
	.datad(Equal6),
	.cin(gnd),
	.combout(\auto_run~0_combout ),
	.cout());
defparam \auto_run~0 .lut_mask = 16'hEFFE;
defparam \auto_run~0 .sum_lutc_input = "datac";

dffeas auto_run(
	.clk(wire_pll7_clk_0),
	.d(\auto_run~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_run~q ),
	.prn(vcc));
defparam auto_run.is_wysiwyg = "true";
defparam auto_run.power_up = "low";

cycloneive_lcell_comb \go~0 (
	.dataa(m0_read),
	.datab(\always0~0_combout ),
	.datac(read_mux_out),
	.datad(\auto_run~q ),
	.cin(gnd),
	.combout(\go~0_combout ),
	.cout());
defparam \go~0 .lut_mask = 16'hFAFC;
defparam \go~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \go~1 (
	.dataa(\go~q ),
	.datab(\go~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\go~1_combout ),
	.cout());
defparam \go~1 .lut_mask = 16'hEEEE;
defparam \go~1 .sum_lutc_input = "datac";

dffeas go(
	.clk(wire_pll7_clk_0),
	.d(\go~1_combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(\ADC_CTRL|currState.doneState~q ),
	.ena(vcc),
	.q(\go~q ),
	.prn(vcc));
defparam go.is_wysiwyg = "true";
defparam go.power_up = "low";

dffeas \values[6][0] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][0]~q ),
	.prn(vcc));
defparam \values[6][0] .is_wysiwyg = "true";
defparam \values[6][0] .power_up = "low";

dffeas \values[5][0] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][0]~q ),
	.prn(vcc));
defparam \values[5][0] .is_wysiwyg = "true";
defparam \values[5][0] .power_up = "low";

dffeas \values[4][0] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][0]~q ),
	.prn(vcc));
defparam \values[4][0] .is_wysiwyg = "true";
defparam \values[4][0] .power_up = "low";

cycloneive_lcell_comb \readdata[0]~0 (
	.dataa(W_alu_result_3),
	.datab(\values[5][0]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][0]~q ),
	.cin(gnd),
	.combout(\readdata[0]~0_combout ),
	.cout());
defparam \readdata[0]~0 .lut_mask = 16'hFFDE;
defparam \readdata[0]~0 .sum_lutc_input = "datac";

dffeas \values[7][0] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][0]~q ),
	.prn(vcc));
defparam \values[7][0] .is_wysiwyg = "true";
defparam \values[7][0] .power_up = "low";

cycloneive_lcell_comb \readdata[0]~1 (
	.dataa(\values[6][0]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[0]~0_combout ),
	.datad(\values[7][0]~q ),
	.cin(gnd),
	.combout(\readdata[0]~1_combout ),
	.cout());
defparam \readdata[0]~1 .lut_mask = 16'hFFBE;
defparam \readdata[0]~1 .sum_lutc_input = "datac";

dffeas \values[2][0] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][0]~q ),
	.prn(vcc));
defparam \values[2][0] .is_wysiwyg = "true";
defparam \values[2][0] .power_up = "low";

dffeas \values[1][0] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][0]~q ),
	.prn(vcc));
defparam \values[1][0] .is_wysiwyg = "true";
defparam \values[1][0] .power_up = "low";

dffeas \values[0][0] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][0]~q ),
	.prn(vcc));
defparam \values[0][0] .is_wysiwyg = "true";
defparam \values[0][0] .power_up = "low";

cycloneive_lcell_comb \readdata[0]~2 (
	.dataa(W_alu_result_3),
	.datab(\values[1][0]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][0]~q ),
	.cin(gnd),
	.combout(\readdata[0]~2_combout ),
	.cout());
defparam \readdata[0]~2 .lut_mask = 16'hFFDE;
defparam \readdata[0]~2 .sum_lutc_input = "datac";

dffeas \values[3][0] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][0]~q ),
	.prn(vcc));
defparam \values[3][0] .is_wysiwyg = "true";
defparam \values[3][0] .power_up = "low";

cycloneive_lcell_comb \readdata[0]~3 (
	.dataa(\values[2][0]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[0]~2_combout ),
	.datad(\values[3][0]~q ),
	.cin(gnd),
	.combout(\readdata[0]~3_combout ),
	.cout());
defparam \readdata[0]~3 .lut_mask = 16'hFFBE;
defparam \readdata[0]~3 .sum_lutc_input = "datac";

dffeas \values[6][1] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][1]~q ),
	.prn(vcc));
defparam \values[6][1] .is_wysiwyg = "true";
defparam \values[6][1] .power_up = "low";

dffeas \values[5][1] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][1]~q ),
	.prn(vcc));
defparam \values[5][1] .is_wysiwyg = "true";
defparam \values[5][1] .power_up = "low";

dffeas \values[4][1] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][1]~q ),
	.prn(vcc));
defparam \values[4][1] .is_wysiwyg = "true";
defparam \values[4][1] .power_up = "low";

cycloneive_lcell_comb \readdata[1]~5 (
	.dataa(W_alu_result_3),
	.datab(\values[5][1]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][1]~q ),
	.cin(gnd),
	.combout(\readdata[1]~5_combout ),
	.cout());
defparam \readdata[1]~5 .lut_mask = 16'hFFDE;
defparam \readdata[1]~5 .sum_lutc_input = "datac";

dffeas \values[7][1] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][1]~q ),
	.prn(vcc));
defparam \values[7][1] .is_wysiwyg = "true";
defparam \values[7][1] .power_up = "low";

cycloneive_lcell_comb \readdata[1]~6 (
	.dataa(\values[6][1]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[1]~5_combout ),
	.datad(\values[7][1]~q ),
	.cin(gnd),
	.combout(\readdata[1]~6_combout ),
	.cout());
defparam \readdata[1]~6 .lut_mask = 16'hFFBE;
defparam \readdata[1]~6 .sum_lutc_input = "datac";

dffeas \values[2][1] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][1]~q ),
	.prn(vcc));
defparam \values[2][1] .is_wysiwyg = "true";
defparam \values[2][1] .power_up = "low";

dffeas \values[1][1] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][1]~q ),
	.prn(vcc));
defparam \values[1][1] .is_wysiwyg = "true";
defparam \values[1][1] .power_up = "low";

dffeas \values[0][1] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][1]~q ),
	.prn(vcc));
defparam \values[0][1] .is_wysiwyg = "true";
defparam \values[0][1] .power_up = "low";

cycloneive_lcell_comb \readdata[1]~7 (
	.dataa(W_alu_result_3),
	.datab(\values[1][1]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][1]~q ),
	.cin(gnd),
	.combout(\readdata[1]~7_combout ),
	.cout());
defparam \readdata[1]~7 .lut_mask = 16'hFFDE;
defparam \readdata[1]~7 .sum_lutc_input = "datac";

dffeas \values[3][1] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][1]~q ),
	.prn(vcc));
defparam \values[3][1] .is_wysiwyg = "true";
defparam \values[3][1] .power_up = "low";

cycloneive_lcell_comb \readdata[1]~8 (
	.dataa(\values[2][1]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[1]~7_combout ),
	.datad(\values[3][1]~q ),
	.cin(gnd),
	.combout(\readdata[1]~8_combout ),
	.cout());
defparam \readdata[1]~8 .lut_mask = 16'hFFBE;
defparam \readdata[1]~8 .sum_lutc_input = "datac";

dffeas \values[6][2] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][2]~q ),
	.prn(vcc));
defparam \values[6][2] .is_wysiwyg = "true";
defparam \values[6][2] .power_up = "low";

dffeas \values[5][2] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][2]~q ),
	.prn(vcc));
defparam \values[5][2] .is_wysiwyg = "true";
defparam \values[5][2] .power_up = "low";

dffeas \values[4][2] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][2]~q ),
	.prn(vcc));
defparam \values[4][2] .is_wysiwyg = "true";
defparam \values[4][2] .power_up = "low";

cycloneive_lcell_comb \readdata[2]~10 (
	.dataa(W_alu_result_3),
	.datab(\values[5][2]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][2]~q ),
	.cin(gnd),
	.combout(\readdata[2]~10_combout ),
	.cout());
defparam \readdata[2]~10 .lut_mask = 16'hFFDE;
defparam \readdata[2]~10 .sum_lutc_input = "datac";

dffeas \values[7][2] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][2]~q ),
	.prn(vcc));
defparam \values[7][2] .is_wysiwyg = "true";
defparam \values[7][2] .power_up = "low";

cycloneive_lcell_comb \readdata[2]~11 (
	.dataa(\values[6][2]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[2]~10_combout ),
	.datad(\values[7][2]~q ),
	.cin(gnd),
	.combout(\readdata[2]~11_combout ),
	.cout());
defparam \readdata[2]~11 .lut_mask = 16'hFFBE;
defparam \readdata[2]~11 .sum_lutc_input = "datac";

dffeas \values[2][2] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][2]~q ),
	.prn(vcc));
defparam \values[2][2] .is_wysiwyg = "true";
defparam \values[2][2] .power_up = "low";

dffeas \values[1][2] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][2]~q ),
	.prn(vcc));
defparam \values[1][2] .is_wysiwyg = "true";
defparam \values[1][2] .power_up = "low";

dffeas \values[0][2] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][2]~q ),
	.prn(vcc));
defparam \values[0][2] .is_wysiwyg = "true";
defparam \values[0][2] .power_up = "low";

cycloneive_lcell_comb \readdata[2]~12 (
	.dataa(W_alu_result_3),
	.datab(\values[1][2]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][2]~q ),
	.cin(gnd),
	.combout(\readdata[2]~12_combout ),
	.cout());
defparam \readdata[2]~12 .lut_mask = 16'hFFDE;
defparam \readdata[2]~12 .sum_lutc_input = "datac";

dffeas \values[3][2] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][2]~q ),
	.prn(vcc));
defparam \values[3][2] .is_wysiwyg = "true";
defparam \values[3][2] .power_up = "low";

cycloneive_lcell_comb \readdata[2]~13 (
	.dataa(\values[2][2]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[2]~12_combout ),
	.datad(\values[3][2]~q ),
	.cin(gnd),
	.combout(\readdata[2]~13_combout ),
	.cout());
defparam \readdata[2]~13 .lut_mask = 16'hFFBE;
defparam \readdata[2]~13 .sum_lutc_input = "datac";

dffeas \values[6][3] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][3]~q ),
	.prn(vcc));
defparam \values[6][3] .is_wysiwyg = "true";
defparam \values[6][3] .power_up = "low";

dffeas \values[5][3] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][3]~q ),
	.prn(vcc));
defparam \values[5][3] .is_wysiwyg = "true";
defparam \values[5][3] .power_up = "low";

dffeas \values[4][3] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][3]~q ),
	.prn(vcc));
defparam \values[4][3] .is_wysiwyg = "true";
defparam \values[4][3] .power_up = "low";

cycloneive_lcell_comb \readdata[3]~15 (
	.dataa(W_alu_result_3),
	.datab(\values[5][3]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][3]~q ),
	.cin(gnd),
	.combout(\readdata[3]~15_combout ),
	.cout());
defparam \readdata[3]~15 .lut_mask = 16'hFFDE;
defparam \readdata[3]~15 .sum_lutc_input = "datac";

dffeas \values[7][3] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][3]~q ),
	.prn(vcc));
defparam \values[7][3] .is_wysiwyg = "true";
defparam \values[7][3] .power_up = "low";

cycloneive_lcell_comb \readdata[3]~16 (
	.dataa(\values[6][3]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[3]~15_combout ),
	.datad(\values[7][3]~q ),
	.cin(gnd),
	.combout(\readdata[3]~16_combout ),
	.cout());
defparam \readdata[3]~16 .lut_mask = 16'hFFBE;
defparam \readdata[3]~16 .sum_lutc_input = "datac";

dffeas \values[2][3] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][3]~q ),
	.prn(vcc));
defparam \values[2][3] .is_wysiwyg = "true";
defparam \values[2][3] .power_up = "low";

dffeas \values[1][3] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][3]~q ),
	.prn(vcc));
defparam \values[1][3] .is_wysiwyg = "true";
defparam \values[1][3] .power_up = "low";

dffeas \values[0][3] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][3]~q ),
	.prn(vcc));
defparam \values[0][3] .is_wysiwyg = "true";
defparam \values[0][3] .power_up = "low";

cycloneive_lcell_comb \readdata[3]~17 (
	.dataa(W_alu_result_3),
	.datab(\values[1][3]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][3]~q ),
	.cin(gnd),
	.combout(\readdata[3]~17_combout ),
	.cout());
defparam \readdata[3]~17 .lut_mask = 16'hFFDE;
defparam \readdata[3]~17 .sum_lutc_input = "datac";

dffeas \values[3][3] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][3]~q ),
	.prn(vcc));
defparam \values[3][3] .is_wysiwyg = "true";
defparam \values[3][3] .power_up = "low";

cycloneive_lcell_comb \readdata[3]~18 (
	.dataa(\values[2][3]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[3]~17_combout ),
	.datad(\values[3][3]~q ),
	.cin(gnd),
	.combout(\readdata[3]~18_combout ),
	.cout());
defparam \readdata[3]~18 .lut_mask = 16'hFFBE;
defparam \readdata[3]~18 .sum_lutc_input = "datac";

dffeas \values[6][4] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][4]~q ),
	.prn(vcc));
defparam \values[6][4] .is_wysiwyg = "true";
defparam \values[6][4] .power_up = "low";

dffeas \values[5][4] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][4]~q ),
	.prn(vcc));
defparam \values[5][4] .is_wysiwyg = "true";
defparam \values[5][4] .power_up = "low";

dffeas \values[4][4] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][4]~q ),
	.prn(vcc));
defparam \values[4][4] .is_wysiwyg = "true";
defparam \values[4][4] .power_up = "low";

cycloneive_lcell_comb \readdata[4]~20 (
	.dataa(W_alu_result_3),
	.datab(\values[5][4]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][4]~q ),
	.cin(gnd),
	.combout(\readdata[4]~20_combout ),
	.cout());
defparam \readdata[4]~20 .lut_mask = 16'hFFDE;
defparam \readdata[4]~20 .sum_lutc_input = "datac";

dffeas \values[7][4] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][4]~q ),
	.prn(vcc));
defparam \values[7][4] .is_wysiwyg = "true";
defparam \values[7][4] .power_up = "low";

cycloneive_lcell_comb \readdata[4]~21 (
	.dataa(\values[6][4]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[4]~20_combout ),
	.datad(\values[7][4]~q ),
	.cin(gnd),
	.combout(\readdata[4]~21_combout ),
	.cout());
defparam \readdata[4]~21 .lut_mask = 16'hFFBE;
defparam \readdata[4]~21 .sum_lutc_input = "datac";

dffeas \values[2][4] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][4]~q ),
	.prn(vcc));
defparam \values[2][4] .is_wysiwyg = "true";
defparam \values[2][4] .power_up = "low";

dffeas \values[1][4] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][4]~q ),
	.prn(vcc));
defparam \values[1][4] .is_wysiwyg = "true";
defparam \values[1][4] .power_up = "low";

dffeas \values[0][4] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][4]~q ),
	.prn(vcc));
defparam \values[0][4] .is_wysiwyg = "true";
defparam \values[0][4] .power_up = "low";

cycloneive_lcell_comb \readdata[4]~22 (
	.dataa(W_alu_result_3),
	.datab(\values[1][4]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][4]~q ),
	.cin(gnd),
	.combout(\readdata[4]~22_combout ),
	.cout());
defparam \readdata[4]~22 .lut_mask = 16'hFFDE;
defparam \readdata[4]~22 .sum_lutc_input = "datac";

dffeas \values[3][4] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][4]~q ),
	.prn(vcc));
defparam \values[3][4] .is_wysiwyg = "true";
defparam \values[3][4] .power_up = "low";

cycloneive_lcell_comb \readdata[4]~23 (
	.dataa(\values[2][4]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[4]~22_combout ),
	.datad(\values[3][4]~q ),
	.cin(gnd),
	.combout(\readdata[4]~23_combout ),
	.cout());
defparam \readdata[4]~23 .lut_mask = 16'hFFBE;
defparam \readdata[4]~23 .sum_lutc_input = "datac";

dffeas \values[6][5] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][5]~q ),
	.prn(vcc));
defparam \values[6][5] .is_wysiwyg = "true";
defparam \values[6][5] .power_up = "low";

dffeas \values[5][5] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][5]~q ),
	.prn(vcc));
defparam \values[5][5] .is_wysiwyg = "true";
defparam \values[5][5] .power_up = "low";

dffeas \values[4][5] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][5]~q ),
	.prn(vcc));
defparam \values[4][5] .is_wysiwyg = "true";
defparam \values[4][5] .power_up = "low";

cycloneive_lcell_comb \readdata[5]~25 (
	.dataa(W_alu_result_3),
	.datab(\values[5][5]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][5]~q ),
	.cin(gnd),
	.combout(\readdata[5]~25_combout ),
	.cout());
defparam \readdata[5]~25 .lut_mask = 16'hFFDE;
defparam \readdata[5]~25 .sum_lutc_input = "datac";

dffeas \values[7][5] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][5]~q ),
	.prn(vcc));
defparam \values[7][5] .is_wysiwyg = "true";
defparam \values[7][5] .power_up = "low";

cycloneive_lcell_comb \readdata[5]~26 (
	.dataa(\values[6][5]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[5]~25_combout ),
	.datad(\values[7][5]~q ),
	.cin(gnd),
	.combout(\readdata[5]~26_combout ),
	.cout());
defparam \readdata[5]~26 .lut_mask = 16'hFFBE;
defparam \readdata[5]~26 .sum_lutc_input = "datac";

dffeas \values[2][5] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][5]~q ),
	.prn(vcc));
defparam \values[2][5] .is_wysiwyg = "true";
defparam \values[2][5] .power_up = "low";

dffeas \values[1][5] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][5]~q ),
	.prn(vcc));
defparam \values[1][5] .is_wysiwyg = "true";
defparam \values[1][5] .power_up = "low";

dffeas \values[0][5] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][5]~q ),
	.prn(vcc));
defparam \values[0][5] .is_wysiwyg = "true";
defparam \values[0][5] .power_up = "low";

cycloneive_lcell_comb \readdata[5]~27 (
	.dataa(W_alu_result_3),
	.datab(\values[1][5]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][5]~q ),
	.cin(gnd),
	.combout(\readdata[5]~27_combout ),
	.cout());
defparam \readdata[5]~27 .lut_mask = 16'hFFDE;
defparam \readdata[5]~27 .sum_lutc_input = "datac";

dffeas \values[3][5] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][5]~q ),
	.prn(vcc));
defparam \values[3][5] .is_wysiwyg = "true";
defparam \values[3][5] .power_up = "low";

cycloneive_lcell_comb \readdata[5]~28 (
	.dataa(\values[2][5]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[5]~27_combout ),
	.datad(\values[3][5]~q ),
	.cin(gnd),
	.combout(\readdata[5]~28_combout ),
	.cout());
defparam \readdata[5]~28 .lut_mask = 16'hFFBE;
defparam \readdata[5]~28 .sum_lutc_input = "datac";

dffeas \values[6][6] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][6]~q ),
	.prn(vcc));
defparam \values[6][6] .is_wysiwyg = "true";
defparam \values[6][6] .power_up = "low";

dffeas \values[5][6] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][6]~q ),
	.prn(vcc));
defparam \values[5][6] .is_wysiwyg = "true";
defparam \values[5][6] .power_up = "low";

dffeas \values[4][6] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][6]~q ),
	.prn(vcc));
defparam \values[4][6] .is_wysiwyg = "true";
defparam \values[4][6] .power_up = "low";

cycloneive_lcell_comb \readdata[6]~30 (
	.dataa(W_alu_result_3),
	.datab(\values[5][6]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][6]~q ),
	.cin(gnd),
	.combout(\readdata[6]~30_combout ),
	.cout());
defparam \readdata[6]~30 .lut_mask = 16'hFFDE;
defparam \readdata[6]~30 .sum_lutc_input = "datac";

dffeas \values[7][6] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][6]~q ),
	.prn(vcc));
defparam \values[7][6] .is_wysiwyg = "true";
defparam \values[7][6] .power_up = "low";

cycloneive_lcell_comb \readdata[6]~31 (
	.dataa(\values[6][6]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[6]~30_combout ),
	.datad(\values[7][6]~q ),
	.cin(gnd),
	.combout(\readdata[6]~31_combout ),
	.cout());
defparam \readdata[6]~31 .lut_mask = 16'hFFBE;
defparam \readdata[6]~31 .sum_lutc_input = "datac";

dffeas \values[2][6] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][6]~q ),
	.prn(vcc));
defparam \values[2][6] .is_wysiwyg = "true";
defparam \values[2][6] .power_up = "low";

dffeas \values[1][6] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][6]~q ),
	.prn(vcc));
defparam \values[1][6] .is_wysiwyg = "true";
defparam \values[1][6] .power_up = "low";

dffeas \values[0][6] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][6]~q ),
	.prn(vcc));
defparam \values[0][6] .is_wysiwyg = "true";
defparam \values[0][6] .power_up = "low";

cycloneive_lcell_comb \readdata[6]~32 (
	.dataa(W_alu_result_3),
	.datab(\values[1][6]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][6]~q ),
	.cin(gnd),
	.combout(\readdata[6]~32_combout ),
	.cout());
defparam \readdata[6]~32 .lut_mask = 16'hFFDE;
defparam \readdata[6]~32 .sum_lutc_input = "datac";

dffeas \values[3][6] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][6]~q ),
	.prn(vcc));
defparam \values[3][6] .is_wysiwyg = "true";
defparam \values[3][6] .power_up = "low";

cycloneive_lcell_comb \readdata[6]~33 (
	.dataa(\values[2][6]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[6]~32_combout ),
	.datad(\values[3][6]~q ),
	.cin(gnd),
	.combout(\readdata[6]~33_combout ),
	.cout());
defparam \readdata[6]~33 .lut_mask = 16'hFFBE;
defparam \readdata[6]~33 .sum_lutc_input = "datac";

dffeas \values[6][7] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][7]~q ),
	.prn(vcc));
defparam \values[6][7] .is_wysiwyg = "true";
defparam \values[6][7] .power_up = "low";

dffeas \values[5][7] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][7]~q ),
	.prn(vcc));
defparam \values[5][7] .is_wysiwyg = "true";
defparam \values[5][7] .power_up = "low";

dffeas \values[4][7] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][7]~q ),
	.prn(vcc));
defparam \values[4][7] .is_wysiwyg = "true";
defparam \values[4][7] .power_up = "low";

cycloneive_lcell_comb \readdata[7]~35 (
	.dataa(W_alu_result_3),
	.datab(\values[5][7]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][7]~q ),
	.cin(gnd),
	.combout(\readdata[7]~35_combout ),
	.cout());
defparam \readdata[7]~35 .lut_mask = 16'hFFDE;
defparam \readdata[7]~35 .sum_lutc_input = "datac";

dffeas \values[7][7] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][7]~q ),
	.prn(vcc));
defparam \values[7][7] .is_wysiwyg = "true";
defparam \values[7][7] .power_up = "low";

cycloneive_lcell_comb \readdata[7]~36 (
	.dataa(\values[6][7]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[7]~35_combout ),
	.datad(\values[7][7]~q ),
	.cin(gnd),
	.combout(\readdata[7]~36_combout ),
	.cout());
defparam \readdata[7]~36 .lut_mask = 16'hFFBE;
defparam \readdata[7]~36 .sum_lutc_input = "datac";

dffeas \values[2][7] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][7]~q ),
	.prn(vcc));
defparam \values[2][7] .is_wysiwyg = "true";
defparam \values[2][7] .power_up = "low";

dffeas \values[1][7] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][7]~q ),
	.prn(vcc));
defparam \values[1][7] .is_wysiwyg = "true";
defparam \values[1][7] .power_up = "low";

dffeas \values[0][7] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][7]~q ),
	.prn(vcc));
defparam \values[0][7] .is_wysiwyg = "true";
defparam \values[0][7] .power_up = "low";

cycloneive_lcell_comb \readdata[7]~37 (
	.dataa(W_alu_result_3),
	.datab(\values[1][7]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][7]~q ),
	.cin(gnd),
	.combout(\readdata[7]~37_combout ),
	.cout());
defparam \readdata[7]~37 .lut_mask = 16'hFFDE;
defparam \readdata[7]~37 .sum_lutc_input = "datac";

dffeas \values[3][7] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][7]~q ),
	.prn(vcc));
defparam \values[3][7] .is_wysiwyg = "true";
defparam \values[3][7] .power_up = "low";

cycloneive_lcell_comb \readdata[7]~38 (
	.dataa(\values[2][7]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[7]~37_combout ),
	.datad(\values[3][7]~q ),
	.cin(gnd),
	.combout(\readdata[7]~38_combout ),
	.cout());
defparam \readdata[7]~38 .lut_mask = 16'hFFBE;
defparam \readdata[7]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(\auto_run~q ),
	.datab(write),
	.datac(Equal3),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hFEFF;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~0 (
	.dataa(W_alu_result_2),
	.datab(W_alu_result_3),
	.datac(W_alu_result_4),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
defparam \Decoder0~0 .lut_mask = 16'hFFFB;
defparam \Decoder0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh~0 (
	.dataa(\refresh[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\refresh~0_combout ),
	.cout());
defparam \refresh~0 .lut_mask = 16'hAAFF;
defparam \refresh~0 .sum_lutc_input = "datac";

dffeas \refresh[5] (
	.clk(wire_pll7_clk_0),
	.d(\refresh~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\ADC_CTRL|currState.doneState~q ),
	.ena(!r_sync_rst),
	.q(\refresh[5]~q ),
	.prn(vcc));
defparam \refresh[5] .is_wysiwyg = "true";
defparam \refresh[5] .power_up = "low";

cycloneive_lcell_comb \Decoder0~1 (
	.dataa(W_alu_result_2),
	.datab(W_alu_result_3),
	.datac(W_alu_result_4),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
defparam \Decoder0~1 .lut_mask = 16'hFFFD;
defparam \Decoder0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh~1 (
	.dataa(\refresh[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~1_combout ),
	.cin(gnd),
	.combout(\refresh~1_combout ),
	.cout());
defparam \refresh~1 .lut_mask = 16'hAAFF;
defparam \refresh~1 .sum_lutc_input = "datac";

dffeas \refresh[6] (
	.clk(wire_pll7_clk_0),
	.d(\refresh~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\ADC_CTRL|currState.doneState~q ),
	.ena(!r_sync_rst),
	.q(\refresh[6]~q ),
	.prn(vcc));
defparam \refresh[6] .is_wysiwyg = "true";
defparam \refresh[6] .power_up = "low";

cycloneive_lcell_comb \Decoder0~2 (
	.dataa(W_alu_result_2),
	.datab(W_alu_result_3),
	.datac(W_alu_result_4),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
defparam \Decoder0~2 .lut_mask = 16'hFFF7;
defparam \Decoder0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh~2 (
	.dataa(\refresh[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\refresh~2_combout ),
	.cout());
defparam \refresh~2 .lut_mask = 16'hAAFF;
defparam \refresh~2 .sum_lutc_input = "datac";

dffeas \refresh[4] (
	.clk(wire_pll7_clk_0),
	.d(\refresh~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\ADC_CTRL|currState.doneState~q ),
	.ena(!r_sync_rst),
	.q(\refresh[4]~q ),
	.prn(vcc));
defparam \refresh[4] .is_wysiwyg = "true";
defparam \refresh[4] .power_up = "low";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(W_alu_result_2),
	.datab(\refresh[6]~q ),
	.datac(W_alu_result_3),
	.datad(\refresh[4]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~3 (
	.dataa(W_alu_result_2),
	.datab(W_alu_result_3),
	.datac(W_alu_result_4),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~3_combout ),
	.cout());
defparam \Decoder0~3 .lut_mask = 16'hFFFE;
defparam \Decoder0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh~3 (
	.dataa(\refresh[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~3_combout ),
	.cin(gnd),
	.combout(\refresh~3_combout ),
	.cout());
defparam \refresh~3 .lut_mask = 16'hAAFF;
defparam \refresh~3 .sum_lutc_input = "datac";

dffeas \refresh[7] (
	.clk(wire_pll7_clk_0),
	.d(\refresh~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\ADC_CTRL|currState.doneState~q ),
	.ena(!r_sync_rst),
	.q(\refresh[7]~q ),
	.prn(vcc));
defparam \refresh[7] .is_wysiwyg = "true";
defparam \refresh[7] .power_up = "low";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\refresh[5]~q ),
	.datab(W_alu_result_2),
	.datac(\Mux0~0_combout ),
	.datad(\refresh[7]~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~4 (
	.dataa(W_alu_result_2),
	.datab(W_alu_result_3),
	.datac(W_alu_result_4),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~4_combout ),
	.cout());
defparam \Decoder0~4 .lut_mask = 16'hFFDF;
defparam \Decoder0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh~4 (
	.dataa(\refresh[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~4_combout ),
	.cin(gnd),
	.combout(\refresh~4_combout ),
	.cout());
defparam \refresh~4 .lut_mask = 16'hAAFF;
defparam \refresh~4 .sum_lutc_input = "datac";

dffeas \refresh[2] (
	.clk(wire_pll7_clk_0),
	.d(\refresh~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\ADC_CTRL|currState.doneState~q ),
	.ena(!r_sync_rst),
	.q(\refresh[2]~q ),
	.prn(vcc));
defparam \refresh[2] .is_wysiwyg = "true";
defparam \refresh[2] .power_up = "low";

cycloneive_lcell_comb \Decoder0~5 (
	.dataa(W_alu_result_2),
	.datab(W_alu_result_3),
	.datac(W_alu_result_4),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~5_combout ),
	.cout());
defparam \Decoder0~5 .lut_mask = 16'hFFBF;
defparam \Decoder0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh~5 (
	.dataa(\refresh[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\refresh~5_combout ),
	.cout());
defparam \refresh~5 .lut_mask = 16'hAAFF;
defparam \refresh~5 .sum_lutc_input = "datac";

dffeas \refresh[1] (
	.clk(wire_pll7_clk_0),
	.d(\refresh~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\ADC_CTRL|currState.doneState~q ),
	.ena(!r_sync_rst),
	.q(\refresh[1]~q ),
	.prn(vcc));
defparam \refresh[1] .is_wysiwyg = "true";
defparam \refresh[1] .power_up = "low";

cycloneive_lcell_comb \Decoder0~6 (
	.dataa(W_alu_result_2),
	.datab(W_alu_result_3),
	.datac(W_alu_result_4),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~6_combout ),
	.cout());
defparam \Decoder0~6 .lut_mask = 16'hFF7F;
defparam \Decoder0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh~6 (
	.dataa(\refresh[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~6_combout ),
	.cin(gnd),
	.combout(\refresh~6_combout ),
	.cout());
defparam \refresh~6 .lut_mask = 16'hAAFF;
defparam \refresh~6 .sum_lutc_input = "datac";

dffeas \refresh[0] (
	.clk(wire_pll7_clk_0),
	.d(\refresh~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\ADC_CTRL|currState.doneState~q ),
	.ena(!r_sync_rst),
	.q(\refresh[0]~q ),
	.prn(vcc));
defparam \refresh[0] .is_wysiwyg = "true";
defparam \refresh[0] .power_up = "low";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(W_alu_result_3),
	.datab(\refresh[1]~q ),
	.datac(W_alu_result_2),
	.datad(\refresh[0]~q ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hFFDE;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~7 (
	.dataa(W_alu_result_2),
	.datab(W_alu_result_3),
	.datac(W_alu_result_4),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~7_combout ),
	.cout());
defparam \Decoder0~7 .lut_mask = 16'hFFEF;
defparam \Decoder0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh~7 (
	.dataa(\refresh[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\refresh~7_combout ),
	.cout());
defparam \refresh~7 .lut_mask = 16'hAAFF;
defparam \refresh~7 .sum_lutc_input = "datac";

dffeas \refresh[3] (
	.clk(wire_pll7_clk_0),
	.d(\refresh~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\ADC_CTRL|currState.doneState~q ),
	.ena(!r_sync_rst),
	.q(\refresh[3]~q ),
	.prn(vcc));
defparam \refresh[3] .is_wysiwyg = "true";
defparam \refresh[3] .power_up = "low";

cycloneive_lcell_comb \Mux0~3 (
	.dataa(\refresh[2]~q ),
	.datab(W_alu_result_3),
	.datac(\Mux0~2_combout ),
	.datad(\refresh[3]~q ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hFFBE;
defparam \Mux0~3 .sum_lutc_input = "datac";

dffeas \values[6][11] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][11]~q ),
	.prn(vcc));
defparam \values[6][11] .is_wysiwyg = "true";
defparam \values[6][11] .power_up = "low";

dffeas \values[5][11] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][11]~q ),
	.prn(vcc));
defparam \values[5][11] .is_wysiwyg = "true";
defparam \values[5][11] .power_up = "low";

dffeas \values[4][11] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][11]~q ),
	.prn(vcc));
defparam \values[4][11] .is_wysiwyg = "true";
defparam \values[4][11] .power_up = "low";

cycloneive_lcell_comb \readdata[11]~41 (
	.dataa(W_alu_result_3),
	.datab(\values[5][11]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][11]~q ),
	.cin(gnd),
	.combout(\readdata[11]~41_combout ),
	.cout());
defparam \readdata[11]~41 .lut_mask = 16'hFFDE;
defparam \readdata[11]~41 .sum_lutc_input = "datac";

dffeas \values[7][11] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][11]~q ),
	.prn(vcc));
defparam \values[7][11] .is_wysiwyg = "true";
defparam \values[7][11] .power_up = "low";

cycloneive_lcell_comb \readdata[11]~42 (
	.dataa(\values[6][11]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[11]~41_combout ),
	.datad(\values[7][11]~q ),
	.cin(gnd),
	.combout(\readdata[11]~42_combout ),
	.cout());
defparam \readdata[11]~42 .lut_mask = 16'hFFBE;
defparam \readdata[11]~42 .sum_lutc_input = "datac";

dffeas \values[2][11] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][11]~q ),
	.prn(vcc));
defparam \values[2][11] .is_wysiwyg = "true";
defparam \values[2][11] .power_up = "low";

dffeas \values[1][11] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][11]~q ),
	.prn(vcc));
defparam \values[1][11] .is_wysiwyg = "true";
defparam \values[1][11] .power_up = "low";

dffeas \values[0][11] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][11]~q ),
	.prn(vcc));
defparam \values[0][11] .is_wysiwyg = "true";
defparam \values[0][11] .power_up = "low";

cycloneive_lcell_comb \readdata[11]~43 (
	.dataa(W_alu_result_3),
	.datab(\values[1][11]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][11]~q ),
	.cin(gnd),
	.combout(\readdata[11]~43_combout ),
	.cout());
defparam \readdata[11]~43 .lut_mask = 16'hFFDE;
defparam \readdata[11]~43 .sum_lutc_input = "datac";

dffeas \values[3][11] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][11]~q ),
	.prn(vcc));
defparam \values[3][11] .is_wysiwyg = "true";
defparam \values[3][11] .power_up = "low";

cycloneive_lcell_comb \readdata[11]~44 (
	.dataa(\values[2][11]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[11]~43_combout ),
	.datad(\values[3][11]~q ),
	.cin(gnd),
	.combout(\readdata[11]~44_combout ),
	.cout());
defparam \readdata[11]~44 .lut_mask = 16'hFFBE;
defparam \readdata[11]~44 .sum_lutc_input = "datac";

dffeas \values[6][10] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][10]~q ),
	.prn(vcc));
defparam \values[6][10] .is_wysiwyg = "true";
defparam \values[6][10] .power_up = "low";

dffeas \values[5][10] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][10]~q ),
	.prn(vcc));
defparam \values[5][10] .is_wysiwyg = "true";
defparam \values[5][10] .power_up = "low";

dffeas \values[4][10] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][10]~q ),
	.prn(vcc));
defparam \values[4][10] .is_wysiwyg = "true";
defparam \values[4][10] .power_up = "low";

cycloneive_lcell_comb \readdata[10]~46 (
	.dataa(W_alu_result_3),
	.datab(\values[5][10]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][10]~q ),
	.cin(gnd),
	.combout(\readdata[10]~46_combout ),
	.cout());
defparam \readdata[10]~46 .lut_mask = 16'hFFDE;
defparam \readdata[10]~46 .sum_lutc_input = "datac";

dffeas \values[7][10] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][10]~q ),
	.prn(vcc));
defparam \values[7][10] .is_wysiwyg = "true";
defparam \values[7][10] .power_up = "low";

cycloneive_lcell_comb \readdata[10]~47 (
	.dataa(\values[6][10]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[10]~46_combout ),
	.datad(\values[7][10]~q ),
	.cin(gnd),
	.combout(\readdata[10]~47_combout ),
	.cout());
defparam \readdata[10]~47 .lut_mask = 16'hFFBE;
defparam \readdata[10]~47 .sum_lutc_input = "datac";

dffeas \values[2][10] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][10]~q ),
	.prn(vcc));
defparam \values[2][10] .is_wysiwyg = "true";
defparam \values[2][10] .power_up = "low";

dffeas \values[1][10] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][10]~q ),
	.prn(vcc));
defparam \values[1][10] .is_wysiwyg = "true";
defparam \values[1][10] .power_up = "low";

dffeas \values[0][10] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][10]~q ),
	.prn(vcc));
defparam \values[0][10] .is_wysiwyg = "true";
defparam \values[0][10] .power_up = "low";

cycloneive_lcell_comb \readdata[10]~48 (
	.dataa(W_alu_result_3),
	.datab(\values[1][10]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][10]~q ),
	.cin(gnd),
	.combout(\readdata[10]~48_combout ),
	.cout());
defparam \readdata[10]~48 .lut_mask = 16'hFFDE;
defparam \readdata[10]~48 .sum_lutc_input = "datac";

dffeas \values[3][10] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][10]~q ),
	.prn(vcc));
defparam \values[3][10] .is_wysiwyg = "true";
defparam \values[3][10] .power_up = "low";

cycloneive_lcell_comb \readdata[10]~49 (
	.dataa(\values[2][10]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[10]~48_combout ),
	.datad(\values[3][10]~q ),
	.cin(gnd),
	.combout(\readdata[10]~49_combout ),
	.cout());
defparam \readdata[10]~49 .lut_mask = 16'hFFBE;
defparam \readdata[10]~49 .sum_lutc_input = "datac";

dffeas \values[6][9] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][9]~q ),
	.prn(vcc));
defparam \values[6][9] .is_wysiwyg = "true";
defparam \values[6][9] .power_up = "low";

dffeas \values[5][9] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][9]~q ),
	.prn(vcc));
defparam \values[5][9] .is_wysiwyg = "true";
defparam \values[5][9] .power_up = "low";

dffeas \values[4][9] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][9]~q ),
	.prn(vcc));
defparam \values[4][9] .is_wysiwyg = "true";
defparam \values[4][9] .power_up = "low";

cycloneive_lcell_comb \readdata[9]~51 (
	.dataa(W_alu_result_3),
	.datab(\values[5][9]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][9]~q ),
	.cin(gnd),
	.combout(\readdata[9]~51_combout ),
	.cout());
defparam \readdata[9]~51 .lut_mask = 16'hFFDE;
defparam \readdata[9]~51 .sum_lutc_input = "datac";

dffeas \values[7][9] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][9]~q ),
	.prn(vcc));
defparam \values[7][9] .is_wysiwyg = "true";
defparam \values[7][9] .power_up = "low";

cycloneive_lcell_comb \readdata[9]~52 (
	.dataa(\values[6][9]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[9]~51_combout ),
	.datad(\values[7][9]~q ),
	.cin(gnd),
	.combout(\readdata[9]~52_combout ),
	.cout());
defparam \readdata[9]~52 .lut_mask = 16'hFFBE;
defparam \readdata[9]~52 .sum_lutc_input = "datac";

dffeas \values[2][9] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][9]~q ),
	.prn(vcc));
defparam \values[2][9] .is_wysiwyg = "true";
defparam \values[2][9] .power_up = "low";

dffeas \values[1][9] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][9]~q ),
	.prn(vcc));
defparam \values[1][9] .is_wysiwyg = "true";
defparam \values[1][9] .power_up = "low";

dffeas \values[0][9] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][9]~q ),
	.prn(vcc));
defparam \values[0][9] .is_wysiwyg = "true";
defparam \values[0][9] .power_up = "low";

cycloneive_lcell_comb \readdata[9]~53 (
	.dataa(W_alu_result_3),
	.datab(\values[1][9]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][9]~q ),
	.cin(gnd),
	.combout(\readdata[9]~53_combout ),
	.cout());
defparam \readdata[9]~53 .lut_mask = 16'hFFDE;
defparam \readdata[9]~53 .sum_lutc_input = "datac";

dffeas \values[3][9] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][9]~q ),
	.prn(vcc));
defparam \values[3][9] .is_wysiwyg = "true";
defparam \values[3][9] .power_up = "low";

cycloneive_lcell_comb \readdata[9]~54 (
	.dataa(\values[2][9]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[9]~53_combout ),
	.datad(\values[3][9]~q ),
	.cin(gnd),
	.combout(\readdata[9]~54_combout ),
	.cout());
defparam \readdata[9]~54 .lut_mask = 16'hFFBE;
defparam \readdata[9]~54 .sum_lutc_input = "datac";

dffeas \values[6][8] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading6[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[6][8]~q ),
	.prn(vcc));
defparam \values[6][8] .is_wysiwyg = "true";
defparam \values[6][8] .power_up = "low";

dffeas \values[5][8] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading5[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[5][8]~q ),
	.prn(vcc));
defparam \values[5][8] .is_wysiwyg = "true";
defparam \values[5][8] .power_up = "low";

dffeas \values[4][8] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading4[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[4][8]~q ),
	.prn(vcc));
defparam \values[4][8] .is_wysiwyg = "true";
defparam \values[4][8] .power_up = "low";

cycloneive_lcell_comb \readdata[8]~56 (
	.dataa(W_alu_result_3),
	.datab(\values[5][8]~q ),
	.datac(W_alu_result_2),
	.datad(\values[4][8]~q ),
	.cin(gnd),
	.combout(\readdata[8]~56_combout ),
	.cout());
defparam \readdata[8]~56 .lut_mask = 16'hFFDE;
defparam \readdata[8]~56 .sum_lutc_input = "datac";

dffeas \values[7][8] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading7[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[7][8]~q ),
	.prn(vcc));
defparam \values[7][8] .is_wysiwyg = "true";
defparam \values[7][8] .power_up = "low";

cycloneive_lcell_comb \readdata[8]~57 (
	.dataa(\values[6][8]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[8]~56_combout ),
	.datad(\values[7][8]~q ),
	.cin(gnd),
	.combout(\readdata[8]~57_combout ),
	.cout());
defparam \readdata[8]~57 .lut_mask = 16'hFFBE;
defparam \readdata[8]~57 .sum_lutc_input = "datac";

dffeas \values[2][8] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading2[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[2][8]~q ),
	.prn(vcc));
defparam \values[2][8] .is_wysiwyg = "true";
defparam \values[2][8] .power_up = "low";

dffeas \values[1][8] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading1[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[1][8]~q ),
	.prn(vcc));
defparam \values[1][8] .is_wysiwyg = "true";
defparam \values[1][8] .power_up = "low";

dffeas \values[0][8] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading0[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[0][8]~q ),
	.prn(vcc));
defparam \values[0][8] .is_wysiwyg = "true";
defparam \values[0][8] .power_up = "low";

cycloneive_lcell_comb \readdata[8]~58 (
	.dataa(W_alu_result_3),
	.datab(\values[1][8]~q ),
	.datac(W_alu_result_2),
	.datad(\values[0][8]~q ),
	.cin(gnd),
	.combout(\readdata[8]~58_combout ),
	.cout());
defparam \readdata[8]~58 .lut_mask = 16'hFFDE;
defparam \readdata[8]~58 .sum_lutc_input = "datac";

dffeas \values[3][8] (
	.clk(wire_pll7_clk_0),
	.d(\ADC_CTRL|reading3[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ADC_CTRL|currState.doneState~q ),
	.q(\values[3][8]~q ),
	.prn(vcc));
defparam \values[3][8] .is_wysiwyg = "true";
defparam \values[3][8] .power_up = "low";

cycloneive_lcell_comb \readdata[8]~59 (
	.dataa(\values[2][8]~q ),
	.datab(W_alu_result_3),
	.datac(\readdata[8]~58_combout ),
	.datad(\values[3][8]~q ),
	.cin(gnd),
	.combout(\readdata[8]~59_combout ),
	.cout());
defparam \readdata[8]~59 .lut_mask = 16'hFFBE;
defparam \readdata[8]~59 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_avalon_adv_adc (
	clock,
	go,
	sclk1,
	cs_n,
	addr_shift_reg_5,
	r_sync_rst,
	currStatedoneState,
	reading6_0,
	reading5_0,
	reading4_0,
	reading7_0,
	reading2_0,
	reading1_0,
	reading0_0,
	reading3_0,
	reading6_1,
	reading5_1,
	reading4_1,
	reading7_1,
	reading2_1,
	reading1_1,
	reading0_1,
	reading3_1,
	reading6_2,
	reading5_2,
	reading4_2,
	reading7_2,
	reading2_2,
	reading1_2,
	reading0_2,
	reading3_2,
	reading6_3,
	reading5_3,
	reading4_3,
	reading7_3,
	reading2_3,
	reading1_3,
	reading0_3,
	reading3_3,
	reading6_4,
	reading5_4,
	reading4_4,
	reading7_4,
	reading2_4,
	reading1_4,
	reading0_4,
	reading3_4,
	reading6_5,
	reading5_5,
	reading4_5,
	reading7_5,
	reading2_5,
	reading1_5,
	reading0_5,
	reading3_5,
	reading6_6,
	reading5_6,
	reading4_6,
	reading7_6,
	reading2_6,
	reading1_6,
	reading0_6,
	reading3_6,
	reading6_7,
	reading5_7,
	reading4_7,
	reading7_7,
	reading2_7,
	reading1_7,
	reading0_7,
	reading3_7,
	reading6_11,
	reading5_11,
	reading4_11,
	reading7_11,
	reading2_11,
	reading1_11,
	reading0_11,
	reading3_11,
	reading6_10,
	reading5_10,
	reading4_10,
	reading7_10,
	reading2_10,
	reading1_10,
	reading0_10,
	reading3_10,
	reading6_9,
	reading5_9,
	reading4_9,
	reading7_9,
	reading2_9,
	reading1_9,
	reading0_9,
	reading3_9,
	reading6_8,
	reading5_8,
	reading4_8,
	reading7_8,
	reading2_8,
	reading1_8,
	reading0_8,
	reading3_8,
	dout)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	go;
output 	sclk1;
output 	cs_n;
output 	addr_shift_reg_5;
input 	r_sync_rst;
output 	currStatedoneState;
output 	reading6_0;
output 	reading5_0;
output 	reading4_0;
output 	reading7_0;
output 	reading2_0;
output 	reading1_0;
output 	reading0_0;
output 	reading3_0;
output 	reading6_1;
output 	reading5_1;
output 	reading4_1;
output 	reading7_1;
output 	reading2_1;
output 	reading1_1;
output 	reading0_1;
output 	reading3_1;
output 	reading6_2;
output 	reading5_2;
output 	reading4_2;
output 	reading7_2;
output 	reading2_2;
output 	reading1_2;
output 	reading0_2;
output 	reading3_2;
output 	reading6_3;
output 	reading5_3;
output 	reading4_3;
output 	reading7_3;
output 	reading2_3;
output 	reading1_3;
output 	reading0_3;
output 	reading3_3;
output 	reading6_4;
output 	reading5_4;
output 	reading4_4;
output 	reading7_4;
output 	reading2_4;
output 	reading1_4;
output 	reading0_4;
output 	reading3_4;
output 	reading6_5;
output 	reading5_5;
output 	reading4_5;
output 	reading7_5;
output 	reading2_5;
output 	reading1_5;
output 	reading0_5;
output 	reading3_5;
output 	reading6_6;
output 	reading5_6;
output 	reading4_6;
output 	reading7_6;
output 	reading2_6;
output 	reading1_6;
output 	reading0_6;
output 	reading3_6;
output 	reading6_7;
output 	reading5_7;
output 	reading4_7;
output 	reading7_7;
output 	reading2_7;
output 	reading1_7;
output 	reading0_7;
output 	reading3_7;
output 	reading6_11;
output 	reading5_11;
output 	reading4_11;
output 	reading7_11;
output 	reading2_11;
output 	reading1_11;
output 	reading0_11;
output 	reading3_11;
output 	reading6_10;
output 	reading5_10;
output 	reading4_10;
output 	reading7_10;
output 	reading2_10;
output 	reading1_10;
output 	reading0_10;
output 	reading3_10;
output 	reading6_9;
output 	reading5_9;
output 	reading4_9;
output 	reading7_9;
output 	reading2_9;
output 	reading1_9;
output 	reading0_9;
output 	reading3_9;
output 	reading6_8;
output 	reading5_8;
output 	reading4_8;
output 	reading7_8;
output 	reading2_8;
output 	reading1_8;
output 	reading0_8;
output 	reading3_8;
input 	dout;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add3~0_combout ;
wire \currState.resetState~q ;
wire \Selector0~0_combout ;
wire \currState.waitState~q ;
wire \Selector1~0_combout ;
wire \next_addr[0]~0_combout ;
wire \next_addr[0]~q ;
wire \Add5~0_combout ;
wire \address~3_combout ;
wire \address[0]~1_combout ;
wire \address[0]~q ;
wire \Add5~2_combout ;
wire \next_addr[1]~q ;
wire \address~2_combout ;
wire \address[1]~q ;
wire \Add5~1_combout ;
wire \next_addr[2]~q ;
wire \address~0_combout ;
wire \address[2]~q ;
wire \Selector1~1_combout ;
wire \sclk_counter~2_combout ;
wire \sclk_counter~5_combout ;
wire \Equal1~1_combout ;
wire \sclk_counter[2]~3_combout ;
wire \sclk_counter[0]~q ;
wire \sclk_counter~6_combout ;
wire \sclk_counter[1]~q ;
wire \sclk_counter~4_combout ;
wire \sclk_counter[2]~q ;
wire \always5~0_combout ;
wire \sclk_counter~7_combout ;
wire \sclk_counter[3]~q ;
wire \Equal1~2_combout ;
wire \Equal1~3_combout ;
wire \always5~1_combout ;
wire \Selector1~2_combout ;
wire \currState.transState~q ;
wire \nextState.pauseState~0_combout ;
wire \currState.pauseState~q ;
wire \counter[7]~12_combout ;
wire \counter[0]~1_combout ;
wire \counter[0]~3_combout ;
wire \counter[0]~_emulated_q ;
wire \counter[0]~2_combout ;
wire \Add3~1 ;
wire \Add3~2_combout ;
wire \counter~11_combout ;
wire \counter[1]~q ;
wire \Add3~3 ;
wire \Add3~4_combout ;
wire \counter~10_combout ;
wire \counter[2]~q ;
wire \Add3~5 ;
wire \Add3~6_combout ;
wire \counter~9_combout ;
wire \counter[3]~q ;
wire \Add3~7 ;
wire \Add3~8_combout ;
wire \counter~8_combout ;
wire \counter[4]~q ;
wire \Add3~9 ;
wire \Add3~10_combout ;
wire \counter~7_combout ;
wire \counter[5]~q ;
wire \Add3~11 ;
wire \Add3~12_combout ;
wire \counter~6_combout ;
wire \counter[6]~q ;
wire \Add3~13 ;
wire \Add3~14_combout ;
wire \counter~5_combout ;
wire \counter[7]~q ;
wire \Equal1~0_combout ;
wire \sclk~0_combout ;
wire \addr_shift_reg~5_combout ;
wire \addr_shift_reg~9_combout ;
wire \addr_shift_reg~10_combout ;
wire \addr_shift_reg[0]~q ;
wire \addr_shift_reg~7_combout ;
wire \addr_shift_reg~8_combout ;
wire \addr_shift_reg[3]~1_combout ;
wire \addr_shift_reg[1]~q ;
wire \addr_shift_reg~4_combout ;
wire \addr_shift_reg~6_combout ;
wire \addr_shift_reg[2]~q ;
wire \addr_shift_reg~3_combout ;
wire \addr_shift_reg[3]~q ;
wire \addr_shift_reg~2_combout ;
wire \addr_shift_reg[4]~q ;
wire \addr_shift_reg~0_combout ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Decoder0~12_combout ;
wire \Decoder0~2_combout ;
wire \Decoder0~3_combout ;
wire \Decoder0~4_combout ;
wire \Decoder0~5_combout ;
wire \Decoder0~6_combout ;
wire \reading7[6]~0_combout ;
wire \Decoder0~7_combout ;
wire \Decoder0~8_combout ;
wire \Decoder0~9_combout ;
wire \Decoder0~10_combout ;
wire \Decoder0~11_combout ;
wire \always7~0_combout ;
wire \shift_reg[0]~q ;
wire \shift_reg[1]~q ;
wire \shift_reg[2]~q ;
wire \shift_reg[3]~q ;
wire \shift_reg[4]~q ;
wire \shift_reg[5]~q ;
wire \shift_reg[6]~q ;
wire \shift_reg[7]~q ;
wire \shift_reg[8]~q ;
wire \shift_reg[9]~q ;
wire \shift_reg[10]~q ;


dffeas sclk(
	.clk(clock),
	.d(\sclk~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sclk1),
	.prn(vcc));
defparam sclk.is_wysiwyg = "true";
defparam sclk.power_up = "low";

cycloneive_lcell_comb \cs_n~2 (
	.dataa(\currState.pauseState~q ),
	.datab(\currState.transState~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(cs_n),
	.cout());
defparam \cs_n~2 .lut_mask = 16'hEEEE;
defparam \cs_n~2 .sum_lutc_input = "datac";

dffeas \addr_shift_reg[5] (
	.clk(clock),
	.d(\addr_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\addr_shift_reg[3]~1_combout ),
	.q(addr_shift_reg_5),
	.prn(vcc));
defparam \addr_shift_reg[5] .is_wysiwyg = "true";
defparam \addr_shift_reg[5] .power_up = "low";

dffeas \currState.doneState (
	.clk(clock),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(currStatedoneState),
	.prn(vcc));
defparam \currState.doneState .is_wysiwyg = "true";
defparam \currState.doneState .power_up = "low";

dffeas \reading6[0] (
	.clk(clock),
	.d(dout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_0),
	.prn(vcc));
defparam \reading6[0] .is_wysiwyg = "true";
defparam \reading6[0] .power_up = "low";

dffeas \reading5[0] (
	.clk(clock),
	.d(dout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_0),
	.prn(vcc));
defparam \reading5[0] .is_wysiwyg = "true";
defparam \reading5[0] .power_up = "low";

dffeas \reading4[0] (
	.clk(clock),
	.d(dout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_0),
	.prn(vcc));
defparam \reading4[0] .is_wysiwyg = "true";
defparam \reading4[0] .power_up = "low";

dffeas \reading7[0] (
	.clk(clock),
	.d(dout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_0),
	.prn(vcc));
defparam \reading7[0] .is_wysiwyg = "true";
defparam \reading7[0] .power_up = "low";

dffeas \reading2[0] (
	.clk(clock),
	.d(dout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_0),
	.prn(vcc));
defparam \reading2[0] .is_wysiwyg = "true";
defparam \reading2[0] .power_up = "low";

dffeas \reading1[0] (
	.clk(clock),
	.d(dout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_0),
	.prn(vcc));
defparam \reading1[0] .is_wysiwyg = "true";
defparam \reading1[0] .power_up = "low";

dffeas \reading0[0] (
	.clk(clock),
	.d(dout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_0),
	.prn(vcc));
defparam \reading0[0] .is_wysiwyg = "true";
defparam \reading0[0] .power_up = "low";

dffeas \reading3[0] (
	.clk(clock),
	.d(dout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_0),
	.prn(vcc));
defparam \reading3[0] .is_wysiwyg = "true";
defparam \reading3[0] .power_up = "low";

dffeas \reading6[1] (
	.clk(clock),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_1),
	.prn(vcc));
defparam \reading6[1] .is_wysiwyg = "true";
defparam \reading6[1] .power_up = "low";

dffeas \reading5[1] (
	.clk(clock),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_1),
	.prn(vcc));
defparam \reading5[1] .is_wysiwyg = "true";
defparam \reading5[1] .power_up = "low";

dffeas \reading4[1] (
	.clk(clock),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_1),
	.prn(vcc));
defparam \reading4[1] .is_wysiwyg = "true";
defparam \reading4[1] .power_up = "low";

dffeas \reading7[1] (
	.clk(clock),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_1),
	.prn(vcc));
defparam \reading7[1] .is_wysiwyg = "true";
defparam \reading7[1] .power_up = "low";

dffeas \reading2[1] (
	.clk(clock),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_1),
	.prn(vcc));
defparam \reading2[1] .is_wysiwyg = "true";
defparam \reading2[1] .power_up = "low";

dffeas \reading1[1] (
	.clk(clock),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_1),
	.prn(vcc));
defparam \reading1[1] .is_wysiwyg = "true";
defparam \reading1[1] .power_up = "low";

dffeas \reading0[1] (
	.clk(clock),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_1),
	.prn(vcc));
defparam \reading0[1] .is_wysiwyg = "true";
defparam \reading0[1] .power_up = "low";

dffeas \reading3[1] (
	.clk(clock),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_1),
	.prn(vcc));
defparam \reading3[1] .is_wysiwyg = "true";
defparam \reading3[1] .power_up = "low";

dffeas \reading6[2] (
	.clk(clock),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_2),
	.prn(vcc));
defparam \reading6[2] .is_wysiwyg = "true";
defparam \reading6[2] .power_up = "low";

dffeas \reading5[2] (
	.clk(clock),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_2),
	.prn(vcc));
defparam \reading5[2] .is_wysiwyg = "true";
defparam \reading5[2] .power_up = "low";

dffeas \reading4[2] (
	.clk(clock),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_2),
	.prn(vcc));
defparam \reading4[2] .is_wysiwyg = "true";
defparam \reading4[2] .power_up = "low";

dffeas \reading7[2] (
	.clk(clock),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_2),
	.prn(vcc));
defparam \reading7[2] .is_wysiwyg = "true";
defparam \reading7[2] .power_up = "low";

dffeas \reading2[2] (
	.clk(clock),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_2),
	.prn(vcc));
defparam \reading2[2] .is_wysiwyg = "true";
defparam \reading2[2] .power_up = "low";

dffeas \reading1[2] (
	.clk(clock),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_2),
	.prn(vcc));
defparam \reading1[2] .is_wysiwyg = "true";
defparam \reading1[2] .power_up = "low";

dffeas \reading0[2] (
	.clk(clock),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_2),
	.prn(vcc));
defparam \reading0[2] .is_wysiwyg = "true";
defparam \reading0[2] .power_up = "low";

dffeas \reading3[2] (
	.clk(clock),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_2),
	.prn(vcc));
defparam \reading3[2] .is_wysiwyg = "true";
defparam \reading3[2] .power_up = "low";

dffeas \reading6[3] (
	.clk(clock),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_3),
	.prn(vcc));
defparam \reading6[3] .is_wysiwyg = "true";
defparam \reading6[3] .power_up = "low";

dffeas \reading5[3] (
	.clk(clock),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_3),
	.prn(vcc));
defparam \reading5[3] .is_wysiwyg = "true";
defparam \reading5[3] .power_up = "low";

dffeas \reading4[3] (
	.clk(clock),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_3),
	.prn(vcc));
defparam \reading4[3] .is_wysiwyg = "true";
defparam \reading4[3] .power_up = "low";

dffeas \reading7[3] (
	.clk(clock),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_3),
	.prn(vcc));
defparam \reading7[3] .is_wysiwyg = "true";
defparam \reading7[3] .power_up = "low";

dffeas \reading2[3] (
	.clk(clock),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_3),
	.prn(vcc));
defparam \reading2[3] .is_wysiwyg = "true";
defparam \reading2[3] .power_up = "low";

dffeas \reading1[3] (
	.clk(clock),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_3),
	.prn(vcc));
defparam \reading1[3] .is_wysiwyg = "true";
defparam \reading1[3] .power_up = "low";

dffeas \reading0[3] (
	.clk(clock),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_3),
	.prn(vcc));
defparam \reading0[3] .is_wysiwyg = "true";
defparam \reading0[3] .power_up = "low";

dffeas \reading3[3] (
	.clk(clock),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_3),
	.prn(vcc));
defparam \reading3[3] .is_wysiwyg = "true";
defparam \reading3[3] .power_up = "low";

dffeas \reading6[4] (
	.clk(clock),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_4),
	.prn(vcc));
defparam \reading6[4] .is_wysiwyg = "true";
defparam \reading6[4] .power_up = "low";

dffeas \reading5[4] (
	.clk(clock),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_4),
	.prn(vcc));
defparam \reading5[4] .is_wysiwyg = "true";
defparam \reading5[4] .power_up = "low";

dffeas \reading4[4] (
	.clk(clock),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_4),
	.prn(vcc));
defparam \reading4[4] .is_wysiwyg = "true";
defparam \reading4[4] .power_up = "low";

dffeas \reading7[4] (
	.clk(clock),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_4),
	.prn(vcc));
defparam \reading7[4] .is_wysiwyg = "true";
defparam \reading7[4] .power_up = "low";

dffeas \reading2[4] (
	.clk(clock),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_4),
	.prn(vcc));
defparam \reading2[4] .is_wysiwyg = "true";
defparam \reading2[4] .power_up = "low";

dffeas \reading1[4] (
	.clk(clock),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_4),
	.prn(vcc));
defparam \reading1[4] .is_wysiwyg = "true";
defparam \reading1[4] .power_up = "low";

dffeas \reading0[4] (
	.clk(clock),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_4),
	.prn(vcc));
defparam \reading0[4] .is_wysiwyg = "true";
defparam \reading0[4] .power_up = "low";

dffeas \reading3[4] (
	.clk(clock),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_4),
	.prn(vcc));
defparam \reading3[4] .is_wysiwyg = "true";
defparam \reading3[4] .power_up = "low";

dffeas \reading6[5] (
	.clk(clock),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_5),
	.prn(vcc));
defparam \reading6[5] .is_wysiwyg = "true";
defparam \reading6[5] .power_up = "low";

dffeas \reading5[5] (
	.clk(clock),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_5),
	.prn(vcc));
defparam \reading5[5] .is_wysiwyg = "true";
defparam \reading5[5] .power_up = "low";

dffeas \reading4[5] (
	.clk(clock),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_5),
	.prn(vcc));
defparam \reading4[5] .is_wysiwyg = "true";
defparam \reading4[5] .power_up = "low";

dffeas \reading7[5] (
	.clk(clock),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_5),
	.prn(vcc));
defparam \reading7[5] .is_wysiwyg = "true";
defparam \reading7[5] .power_up = "low";

dffeas \reading2[5] (
	.clk(clock),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_5),
	.prn(vcc));
defparam \reading2[5] .is_wysiwyg = "true";
defparam \reading2[5] .power_up = "low";

dffeas \reading1[5] (
	.clk(clock),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_5),
	.prn(vcc));
defparam \reading1[5] .is_wysiwyg = "true";
defparam \reading1[5] .power_up = "low";

dffeas \reading0[5] (
	.clk(clock),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_5),
	.prn(vcc));
defparam \reading0[5] .is_wysiwyg = "true";
defparam \reading0[5] .power_up = "low";

dffeas \reading3[5] (
	.clk(clock),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_5),
	.prn(vcc));
defparam \reading3[5] .is_wysiwyg = "true";
defparam \reading3[5] .power_up = "low";

dffeas \reading6[6] (
	.clk(clock),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_6),
	.prn(vcc));
defparam \reading6[6] .is_wysiwyg = "true";
defparam \reading6[6] .power_up = "low";

dffeas \reading5[6] (
	.clk(clock),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_6),
	.prn(vcc));
defparam \reading5[6] .is_wysiwyg = "true";
defparam \reading5[6] .power_up = "low";

dffeas \reading4[6] (
	.clk(clock),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_6),
	.prn(vcc));
defparam \reading4[6] .is_wysiwyg = "true";
defparam \reading4[6] .power_up = "low";

dffeas \reading7[6] (
	.clk(clock),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_6),
	.prn(vcc));
defparam \reading7[6] .is_wysiwyg = "true";
defparam \reading7[6] .power_up = "low";

dffeas \reading2[6] (
	.clk(clock),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_6),
	.prn(vcc));
defparam \reading2[6] .is_wysiwyg = "true";
defparam \reading2[6] .power_up = "low";

dffeas \reading1[6] (
	.clk(clock),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_6),
	.prn(vcc));
defparam \reading1[6] .is_wysiwyg = "true";
defparam \reading1[6] .power_up = "low";

dffeas \reading0[6] (
	.clk(clock),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_6),
	.prn(vcc));
defparam \reading0[6] .is_wysiwyg = "true";
defparam \reading0[6] .power_up = "low";

dffeas \reading3[6] (
	.clk(clock),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_6),
	.prn(vcc));
defparam \reading3[6] .is_wysiwyg = "true";
defparam \reading3[6] .power_up = "low";

dffeas \reading6[7] (
	.clk(clock),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_7),
	.prn(vcc));
defparam \reading6[7] .is_wysiwyg = "true";
defparam \reading6[7] .power_up = "low";

dffeas \reading5[7] (
	.clk(clock),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_7),
	.prn(vcc));
defparam \reading5[7] .is_wysiwyg = "true";
defparam \reading5[7] .power_up = "low";

dffeas \reading4[7] (
	.clk(clock),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_7),
	.prn(vcc));
defparam \reading4[7] .is_wysiwyg = "true";
defparam \reading4[7] .power_up = "low";

dffeas \reading7[7] (
	.clk(clock),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_7),
	.prn(vcc));
defparam \reading7[7] .is_wysiwyg = "true";
defparam \reading7[7] .power_up = "low";

dffeas \reading2[7] (
	.clk(clock),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_7),
	.prn(vcc));
defparam \reading2[7] .is_wysiwyg = "true";
defparam \reading2[7] .power_up = "low";

dffeas \reading1[7] (
	.clk(clock),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_7),
	.prn(vcc));
defparam \reading1[7] .is_wysiwyg = "true";
defparam \reading1[7] .power_up = "low";

dffeas \reading0[7] (
	.clk(clock),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_7),
	.prn(vcc));
defparam \reading0[7] .is_wysiwyg = "true";
defparam \reading0[7] .power_up = "low";

dffeas \reading3[7] (
	.clk(clock),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_7),
	.prn(vcc));
defparam \reading3[7] .is_wysiwyg = "true";
defparam \reading3[7] .power_up = "low";

dffeas \reading6[11] (
	.clk(clock),
	.d(\shift_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_11),
	.prn(vcc));
defparam \reading6[11] .is_wysiwyg = "true";
defparam \reading6[11] .power_up = "low";

dffeas \reading5[11] (
	.clk(clock),
	.d(\shift_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_11),
	.prn(vcc));
defparam \reading5[11] .is_wysiwyg = "true";
defparam \reading5[11] .power_up = "low";

dffeas \reading4[11] (
	.clk(clock),
	.d(\shift_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_11),
	.prn(vcc));
defparam \reading4[11] .is_wysiwyg = "true";
defparam \reading4[11] .power_up = "low";

dffeas \reading7[11] (
	.clk(clock),
	.d(\shift_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_11),
	.prn(vcc));
defparam \reading7[11] .is_wysiwyg = "true";
defparam \reading7[11] .power_up = "low";

dffeas \reading2[11] (
	.clk(clock),
	.d(\shift_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_11),
	.prn(vcc));
defparam \reading2[11] .is_wysiwyg = "true";
defparam \reading2[11] .power_up = "low";

dffeas \reading1[11] (
	.clk(clock),
	.d(\shift_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_11),
	.prn(vcc));
defparam \reading1[11] .is_wysiwyg = "true";
defparam \reading1[11] .power_up = "low";

dffeas \reading0[11] (
	.clk(clock),
	.d(\shift_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_11),
	.prn(vcc));
defparam \reading0[11] .is_wysiwyg = "true";
defparam \reading0[11] .power_up = "low";

dffeas \reading3[11] (
	.clk(clock),
	.d(\shift_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_11),
	.prn(vcc));
defparam \reading3[11] .is_wysiwyg = "true";
defparam \reading3[11] .power_up = "low";

dffeas \reading6[10] (
	.clk(clock),
	.d(\shift_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_10),
	.prn(vcc));
defparam \reading6[10] .is_wysiwyg = "true";
defparam \reading6[10] .power_up = "low";

dffeas \reading5[10] (
	.clk(clock),
	.d(\shift_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_10),
	.prn(vcc));
defparam \reading5[10] .is_wysiwyg = "true";
defparam \reading5[10] .power_up = "low";

dffeas \reading4[10] (
	.clk(clock),
	.d(\shift_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_10),
	.prn(vcc));
defparam \reading4[10] .is_wysiwyg = "true";
defparam \reading4[10] .power_up = "low";

dffeas \reading7[10] (
	.clk(clock),
	.d(\shift_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_10),
	.prn(vcc));
defparam \reading7[10] .is_wysiwyg = "true";
defparam \reading7[10] .power_up = "low";

dffeas \reading2[10] (
	.clk(clock),
	.d(\shift_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_10),
	.prn(vcc));
defparam \reading2[10] .is_wysiwyg = "true";
defparam \reading2[10] .power_up = "low";

dffeas \reading1[10] (
	.clk(clock),
	.d(\shift_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_10),
	.prn(vcc));
defparam \reading1[10] .is_wysiwyg = "true";
defparam \reading1[10] .power_up = "low";

dffeas \reading0[10] (
	.clk(clock),
	.d(\shift_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_10),
	.prn(vcc));
defparam \reading0[10] .is_wysiwyg = "true";
defparam \reading0[10] .power_up = "low";

dffeas \reading3[10] (
	.clk(clock),
	.d(\shift_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_10),
	.prn(vcc));
defparam \reading3[10] .is_wysiwyg = "true";
defparam \reading3[10] .power_up = "low";

dffeas \reading6[9] (
	.clk(clock),
	.d(\shift_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_9),
	.prn(vcc));
defparam \reading6[9] .is_wysiwyg = "true";
defparam \reading6[9] .power_up = "low";

dffeas \reading5[9] (
	.clk(clock),
	.d(\shift_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_9),
	.prn(vcc));
defparam \reading5[9] .is_wysiwyg = "true";
defparam \reading5[9] .power_up = "low";

dffeas \reading4[9] (
	.clk(clock),
	.d(\shift_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_9),
	.prn(vcc));
defparam \reading4[9] .is_wysiwyg = "true";
defparam \reading4[9] .power_up = "low";

dffeas \reading7[9] (
	.clk(clock),
	.d(\shift_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_9),
	.prn(vcc));
defparam \reading7[9] .is_wysiwyg = "true";
defparam \reading7[9] .power_up = "low";

dffeas \reading2[9] (
	.clk(clock),
	.d(\shift_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_9),
	.prn(vcc));
defparam \reading2[9] .is_wysiwyg = "true";
defparam \reading2[9] .power_up = "low";

dffeas \reading1[9] (
	.clk(clock),
	.d(\shift_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_9),
	.prn(vcc));
defparam \reading1[9] .is_wysiwyg = "true";
defparam \reading1[9] .power_up = "low";

dffeas \reading0[9] (
	.clk(clock),
	.d(\shift_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_9),
	.prn(vcc));
defparam \reading0[9] .is_wysiwyg = "true";
defparam \reading0[9] .power_up = "low";

dffeas \reading3[9] (
	.clk(clock),
	.d(\shift_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_9),
	.prn(vcc));
defparam \reading3[9] .is_wysiwyg = "true";
defparam \reading3[9] .power_up = "low";

dffeas \reading6[8] (
	.clk(clock),
	.d(\shift_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.q(reading6_8),
	.prn(vcc));
defparam \reading6[8] .is_wysiwyg = "true";
defparam \reading6[8] .power_up = "low";

dffeas \reading5[8] (
	.clk(clock),
	.d(\shift_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.q(reading5_8),
	.prn(vcc));
defparam \reading5[8] .is_wysiwyg = "true";
defparam \reading5[8] .power_up = "low";

dffeas \reading4[8] (
	.clk(clock),
	.d(\shift_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.q(reading4_8),
	.prn(vcc));
defparam \reading4[8] .is_wysiwyg = "true";
defparam \reading4[8] .power_up = "low";

dffeas \reading7[8] (
	.clk(clock),
	.d(\shift_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\reading7[6]~0_combout ),
	.q(reading7_8),
	.prn(vcc));
defparam \reading7[8] .is_wysiwyg = "true";
defparam \reading7[8] .power_up = "low";

dffeas \reading2[8] (
	.clk(clock),
	.d(\shift_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.q(reading2_8),
	.prn(vcc));
defparam \reading2[8] .is_wysiwyg = "true";
defparam \reading2[8] .power_up = "low";

dffeas \reading1[8] (
	.clk(clock),
	.d(\shift_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.q(reading1_8),
	.prn(vcc));
defparam \reading1[8] .is_wysiwyg = "true";
defparam \reading1[8] .power_up = "low";

dffeas \reading0[8] (
	.clk(clock),
	.d(\shift_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.q(reading0_8),
	.prn(vcc));
defparam \reading0[8] .is_wysiwyg = "true";
defparam \reading0[8] .power_up = "low";

dffeas \reading3[8] (
	.clk(clock),
	.d(\shift_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.q(reading3_8),
	.prn(vcc));
defparam \reading3[8] .is_wysiwyg = "true";
defparam \reading3[8] .power_up = "low";

cycloneive_lcell_comb \Add3~0 (
	.dataa(\counter[0]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout(\Add3~1 ));
defparam \Add3~0 .lut_mask = 16'h55AA;
defparam \Add3~0 .sum_lutc_input = "datac";

dffeas \currState.resetState (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\currState.resetState~q ),
	.prn(vcc));
defparam \currState.resetState .is_wysiwyg = "true";
defparam \currState.resetState .power_up = "low";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\currState.waitState~q ),
	.datab(currStatedoneState),
	.datac(go),
	.datad(\currState.resetState~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEFFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

dffeas \currState.waitState (
	.clk(clock),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\currState.waitState~q ),
	.prn(vcc));
defparam \currState.waitState .is_wysiwyg = "true";
defparam \currState.waitState .power_up = "low";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(go),
	.datab(\currState.waitState~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hEEEE;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_addr[0]~0 (
	.dataa(\address[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_addr[0]~0_combout ),
	.cout());
defparam \next_addr[0]~0 .lut_mask = 16'h5555;
defparam \next_addr[0]~0 .sum_lutc_input = "datac";

dffeas \next_addr[0] (
	.clk(clock),
	.d(\next_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\next_addr[0]~q ),
	.prn(vcc));
defparam \next_addr[0] .is_wysiwyg = "true";
defparam \next_addr[0] .power_up = "low";

cycloneive_lcell_comb \Add5~0 (
	.dataa(\address[1]~q ),
	.datab(\address[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add5~0_combout ),
	.cout());
defparam \Add5~0 .lut_mask = 16'hEEEE;
defparam \Add5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address~3 (
	.dataa(\next_addr[0]~q ),
	.datab(\address[2]~q ),
	.datac(\Add5~0_combout ),
	.datad(\currState.resetState~q ),
	.cin(gnd),
	.combout(\address~3_combout ),
	.cout());
defparam \address~3 .lut_mask = 16'hBFFF;
defparam \address~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address[0]~1 (
	.dataa(\currState.pauseState~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\currState.resetState~q ),
	.cin(gnd),
	.combout(\address[0]~1_combout ),
	.cout());
defparam \address[0]~1 .lut_mask = 16'hAAFF;
defparam \address[0]~1 .sum_lutc_input = "datac";

dffeas \address[0] (
	.clk(clock),
	.d(\address~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[0]~1_combout ),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

cycloneive_lcell_comb \Add5~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\address[1]~q ),
	.datad(\address[0]~q ),
	.cin(gnd),
	.combout(\Add5~2_combout ),
	.cout());
defparam \Add5~2 .lut_mask = 16'h0FF0;
defparam \Add5~2 .sum_lutc_input = "datac";

dffeas \next_addr[1] (
	.clk(clock),
	.d(\Add5~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\next_addr[1]~q ),
	.prn(vcc));
defparam \next_addr[1] .is_wysiwyg = "true";
defparam \next_addr[1] .power_up = "low";

cycloneive_lcell_comb \address~2 (
	.dataa(\currState.resetState~q ),
	.datab(\next_addr[1]~q ),
	.datac(\address[2]~q ),
	.datad(\Add5~0_combout ),
	.cin(gnd),
	.combout(\address~2_combout ),
	.cout());
defparam \address~2 .lut_mask = 16'hEFFF;
defparam \address~2 .sum_lutc_input = "datac";

dffeas \address[1] (
	.clk(clock),
	.d(\address~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[0]~1_combout ),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

cycloneive_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(\address[2]~q ),
	.datac(\address[1]~q ),
	.datad(\address[0]~q ),
	.cin(gnd),
	.combout(\Add5~1_combout ),
	.cout());
defparam \Add5~1 .lut_mask = 16'hC33C;
defparam \Add5~1 .sum_lutc_input = "datac";

dffeas \next_addr[2] (
	.clk(clock),
	.d(\Add5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\next_addr[2]~q ),
	.prn(vcc));
defparam \next_addr[2] .is_wysiwyg = "true";
defparam \next_addr[2] .power_up = "low";

cycloneive_lcell_comb \address~0 (
	.dataa(\currState.resetState~q ),
	.datab(\next_addr[2]~q ),
	.datac(\address[2]~q ),
	.datad(\Add5~0_combout ),
	.cin(gnd),
	.combout(\address~0_combout ),
	.cout());
defparam \address~0 .lut_mask = 16'hEFFF;
defparam \address~0 .sum_lutc_input = "datac";

dffeas \address[2] (
	.clk(clock),
	.d(\address~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[0]~1_combout ),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

cycloneive_lcell_comb \Selector1~1 (
	.dataa(\currState.pauseState~q ),
	.datab(\address[2]~q ),
	.datac(\address[1]~q ),
	.datad(\address[0]~q ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hFFFE;
defparam \Selector1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sclk_counter~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\currState.waitState~q ),
	.datad(currStatedoneState),
	.cin(gnd),
	.combout(\sclk_counter~2_combout ),
	.cout());
defparam \sclk_counter~2 .lut_mask = 16'h0FFF;
defparam \sclk_counter~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sclk_counter~5 (
	.dataa(\sclk_counter[0]~q ),
	.datab(\currState.waitState~q ),
	.datac(currStatedoneState),
	.datad(gnd),
	.cin(gnd),
	.combout(\sclk_counter~5_combout ),
	.cout());
defparam \sclk_counter~5 .lut_mask = 16'h7F7F;
defparam \sclk_counter~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(\counter[0]~2_combout ),
	.datab(\counter[3]~q ),
	.datac(\counter[2]~q ),
	.datad(\counter[1]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hBFFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sclk_counter[2]~3 (
	.dataa(\sclk_counter~2_combout ),
	.datab(\Equal1~0_combout ),
	.datac(\Equal1~1_combout ),
	.datad(sclk1),
	.cin(gnd),
	.combout(\sclk_counter[2]~3_combout ),
	.cout());
defparam \sclk_counter[2]~3 .lut_mask = 16'hFF7F;
defparam \sclk_counter[2]~3 .sum_lutc_input = "datac";

dffeas \sclk_counter[0] (
	.clk(clock),
	.d(\sclk_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sclk_counter[2]~3_combout ),
	.q(\sclk_counter[0]~q ),
	.prn(vcc));
defparam \sclk_counter[0] .is_wysiwyg = "true";
defparam \sclk_counter[0] .power_up = "low";

cycloneive_lcell_comb \sclk_counter~6 (
	.dataa(\sclk_counter[0]~q ),
	.datab(\sclk_counter[1]~q ),
	.datac(\currState.waitState~q ),
	.datad(currStatedoneState),
	.cin(gnd),
	.combout(\sclk_counter~6_combout ),
	.cout());
defparam \sclk_counter~6 .lut_mask = 16'h6FFF;
defparam \sclk_counter~6 .sum_lutc_input = "datac";

dffeas \sclk_counter[1] (
	.clk(clock),
	.d(\sclk_counter~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sclk_counter[2]~3_combout ),
	.q(\sclk_counter[1]~q ),
	.prn(vcc));
defparam \sclk_counter[1] .is_wysiwyg = "true";
defparam \sclk_counter[1] .power_up = "low";

cycloneive_lcell_comb \sclk_counter~4 (
	.dataa(\sclk_counter~2_combout ),
	.datab(\sclk_counter[2]~q ),
	.datac(\sclk_counter[0]~q ),
	.datad(\sclk_counter[1]~q ),
	.cin(gnd),
	.combout(\sclk_counter~4_combout ),
	.cout());
defparam \sclk_counter~4 .lut_mask = 16'hEBBE;
defparam \sclk_counter~4 .sum_lutc_input = "datac";

dffeas \sclk_counter[2] (
	.clk(clock),
	.d(\sclk_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sclk_counter[2]~3_combout ),
	.q(\sclk_counter[2]~q ),
	.prn(vcc));
defparam \sclk_counter[2] .is_wysiwyg = "true";
defparam \sclk_counter[2] .power_up = "low";

cycloneive_lcell_comb \always5~0 (
	.dataa(\sclk_counter[2]~q ),
	.datab(\sclk_counter[0]~q ),
	.datac(\sclk_counter[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'hFEFE;
defparam \always5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sclk_counter~7 (
	.dataa(\currState.waitState~q ),
	.datab(currStatedoneState),
	.datac(\sclk_counter[3]~q ),
	.datad(\always5~0_combout ),
	.cin(gnd),
	.combout(\sclk_counter~7_combout ),
	.cout());
defparam \sclk_counter~7 .lut_mask = 16'h7FF7;
defparam \sclk_counter~7 .sum_lutc_input = "datac";

dffeas \sclk_counter[3] (
	.clk(clock),
	.d(\sclk_counter~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sclk_counter[2]~3_combout ),
	.q(\sclk_counter[3]~q ),
	.prn(vcc));
defparam \sclk_counter[3] .is_wysiwyg = "true";
defparam \sclk_counter[3] .power_up = "low";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(\counter[3]~q ),
	.datab(\counter[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'h7777;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~3 (
	.dataa(\Equal1~0_combout ),
	.datab(\counter[0]~2_combout ),
	.datac(\counter[1]~q ),
	.datad(\Equal1~2_combout ),
	.cin(gnd),
	.combout(\Equal1~3_combout ),
	.cout());
defparam \Equal1~3 .lut_mask = 16'hFFEF;
defparam \Equal1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always5~1 (
	.dataa(sclk1),
	.datab(\sclk_counter[3]~q ),
	.datac(\always5~0_combout ),
	.datad(\Equal1~3_combout ),
	.cin(gnd),
	.combout(\always5~1_combout ),
	.cout());
defparam \always5~1 .lut_mask = 16'hFEFF;
defparam \always5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~2 (
	.dataa(\Selector1~0_combout ),
	.datab(\Selector1~1_combout ),
	.datac(\currState.transState~q ),
	.datad(\always5~1_combout ),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hFEFF;
defparam \Selector1~2 .sum_lutc_input = "datac";

dffeas \currState.transState (
	.clk(clock),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\currState.transState~q ),
	.prn(vcc));
defparam \currState.transState .is_wysiwyg = "true";
defparam \currState.transState .power_up = "low";

cycloneive_lcell_comb \nextState.pauseState~0 (
	.dataa(\currState.transState~q ),
	.datab(\always5~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nextState.pauseState~0_combout ),
	.cout());
defparam \nextState.pauseState~0 .lut_mask = 16'hEEEE;
defparam \nextState.pauseState~0 .sum_lutc_input = "datac";

dffeas \currState.pauseState (
	.clk(clock),
	.d(\nextState.pauseState~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\currState.pauseState~q ),
	.prn(vcc));
defparam \currState.pauseState .is_wysiwyg = "true";
defparam \currState.pauseState .power_up = "low";

cycloneive_lcell_comb \counter[7]~12 (
	.dataa(\currState.pauseState~q ),
	.datab(\currState.transState~q ),
	.datac(\Equal1~0_combout ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\counter[7]~12_combout ),
	.cout());
defparam \counter[7]~12 .lut_mask = 16'hFFFE;
defparam \counter[7]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter[0]~1 (
	.dataa(gnd),
	.datab(sclk1),
	.datac(\counter[0]~1_combout ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\counter[0]~1_combout ),
	.cout());
defparam \counter[0]~1 .lut_mask = 16'hF033;
defparam \counter[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter[0]~3 (
	.dataa(\Add3~0_combout ),
	.datab(\counter[7]~12_combout ),
	.datac(sclk1),
	.datad(\counter[0]~1_combout ),
	.cin(gnd),
	.combout(\counter[0]~3_combout ),
	.cout());
defparam \counter[0]~3 .lut_mask = 16'h6996;
defparam \counter[0]~3 .sum_lutc_input = "datac";

dffeas \counter[0]~_emulated (
	.clk(clock),
	.d(\counter[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter[0]~_emulated_q ),
	.prn(vcc));
defparam \counter[0]~_emulated .is_wysiwyg = "true";
defparam \counter[0]~_emulated .power_up = "low";

cycloneive_lcell_comb \counter[0]~2 (
	.dataa(\counter[0]~_emulated_q ),
	.datab(\counter[0]~1_combout ),
	.datac(r_sync_rst),
	.datad(sclk1),
	.cin(gnd),
	.combout(\counter[0]~2_combout ),
	.cout());
defparam \counter[0]~2 .lut_mask = 16'h96FF;
defparam \counter[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~2 (
	.dataa(\counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~1 ),
	.combout(\Add3~2_combout ),
	.cout(\Add3~3 ));
defparam \Add3~2 .lut_mask = 16'h5AAF;
defparam \Add3~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \counter~11 (
	.dataa(\Add3~2_combout ),
	.datab(\Equal1~0_combout ),
	.datac(\Equal1~1_combout ),
	.datad(cs_n),
	.cin(gnd),
	.combout(\counter~11_combout ),
	.cout());
defparam \counter~11 .lut_mask = 16'hFFFD;
defparam \counter~11 .sum_lutc_input = "datac";

dffeas \counter[1] (
	.clk(clock),
	.d(\counter~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter[1]~q ),
	.prn(vcc));
defparam \counter[1] .is_wysiwyg = "true";
defparam \counter[1] .power_up = "low";

cycloneive_lcell_comb \Add3~4 (
	.dataa(\counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~3 ),
	.combout(\Add3~4_combout ),
	.cout(\Add3~5 ));
defparam \Add3~4 .lut_mask = 16'h5A5F;
defparam \Add3~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \counter~10 (
	.dataa(\Add3~4_combout ),
	.datab(\Equal1~0_combout ),
	.datac(\Equal1~1_combout ),
	.datad(cs_n),
	.cin(gnd),
	.combout(\counter~10_combout ),
	.cout());
defparam \counter~10 .lut_mask = 16'hFFFD;
defparam \counter~10 .sum_lutc_input = "datac";

dffeas \counter[2] (
	.clk(clock),
	.d(\counter~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter[2]~q ),
	.prn(vcc));
defparam \counter[2] .is_wysiwyg = "true";
defparam \counter[2] .power_up = "low";

cycloneive_lcell_comb \Add3~6 (
	.dataa(\counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~5 ),
	.combout(\Add3~6_combout ),
	.cout(\Add3~7 ));
defparam \Add3~6 .lut_mask = 16'h5AAF;
defparam \Add3~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \counter~9 (
	.dataa(\Add3~6_combout ),
	.datab(\Equal1~0_combout ),
	.datac(\Equal1~1_combout ),
	.datad(cs_n),
	.cin(gnd),
	.combout(\counter~9_combout ),
	.cout());
defparam \counter~9 .lut_mask = 16'hFFFD;
defparam \counter~9 .sum_lutc_input = "datac";

dffeas \counter[3] (
	.clk(clock),
	.d(\counter~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter[3]~q ),
	.prn(vcc));
defparam \counter[3] .is_wysiwyg = "true";
defparam \counter[3] .power_up = "low";

cycloneive_lcell_comb \Add3~8 (
	.dataa(\counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~7 ),
	.combout(\Add3~8_combout ),
	.cout(\Add3~9 ));
defparam \Add3~8 .lut_mask = 16'h5AAF;
defparam \Add3~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \counter~8 (
	.dataa(cs_n),
	.datab(\Add3~8_combout ),
	.datac(\Equal1~0_combout ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\counter~8_combout ),
	.cout());
defparam \counter~8 .lut_mask = 16'hFFFE;
defparam \counter~8 .sum_lutc_input = "datac";

dffeas \counter[4] (
	.clk(clock),
	.d(\counter~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter[4]~q ),
	.prn(vcc));
defparam \counter[4] .is_wysiwyg = "true";
defparam \counter[4] .power_up = "low";

cycloneive_lcell_comb \Add3~10 (
	.dataa(\counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~9 ),
	.combout(\Add3~10_combout ),
	.cout(\Add3~11 ));
defparam \Add3~10 .lut_mask = 16'h5A5F;
defparam \Add3~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \counter~7 (
	.dataa(cs_n),
	.datab(\Add3~10_combout ),
	.datac(\Equal1~0_combout ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\counter~7_combout ),
	.cout());
defparam \counter~7 .lut_mask = 16'hFFFE;
defparam \counter~7 .sum_lutc_input = "datac";

dffeas \counter[5] (
	.clk(clock),
	.d(\counter~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter[5]~q ),
	.prn(vcc));
defparam \counter[5] .is_wysiwyg = "true";
defparam \counter[5] .power_up = "low";

cycloneive_lcell_comb \Add3~12 (
	.dataa(\counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~11 ),
	.combout(\Add3~12_combout ),
	.cout(\Add3~13 ));
defparam \Add3~12 .lut_mask = 16'h5AAF;
defparam \Add3~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \counter~6 (
	.dataa(cs_n),
	.datab(\Add3~12_combout ),
	.datac(\Equal1~0_combout ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\counter~6_combout ),
	.cout());
defparam \counter~6 .lut_mask = 16'hFFFE;
defparam \counter~6 .sum_lutc_input = "datac";

dffeas \counter[6] (
	.clk(clock),
	.d(\counter~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter[6]~q ),
	.prn(vcc));
defparam \counter[6] .is_wysiwyg = "true";
defparam \counter[6] .power_up = "low";

cycloneive_lcell_comb \Add3~14 (
	.dataa(\counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add3~13 ),
	.combout(\Add3~14_combout ),
	.cout());
defparam \Add3~14 .lut_mask = 16'h5A5A;
defparam \Add3~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \counter~5 (
	.dataa(cs_n),
	.datab(\Add3~14_combout ),
	.datac(\Equal1~0_combout ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\counter~5_combout ),
	.cout());
defparam \counter~5 .lut_mask = 16'hFFFE;
defparam \counter~5 .sum_lutc_input = "datac";

dffeas \counter[7] (
	.clk(clock),
	.d(\counter~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter[7]~q ),
	.prn(vcc));
defparam \counter[7] .is_wysiwyg = "true";
defparam \counter[7] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\counter[7]~q ),
	.datab(\counter[6]~q ),
	.datac(\counter[5]~q ),
	.datad(\counter[4]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hFFFE;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sclk~0 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(sclk1),
	.datad(cs_n),
	.cin(gnd),
	.combout(\sclk~0_combout ),
	.cout());
defparam \sclk~0 .lut_mask = 16'hFF96;
defparam \sclk~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_shift_reg~5 (
	.dataa(\currState.pauseState~q ),
	.datab(\address[2]~q ),
	.datac(\address[1]~q ),
	.datad(\address[0]~q ),
	.cin(gnd),
	.combout(\addr_shift_reg~5_combout ),
	.cout());
defparam \addr_shift_reg~5 .lut_mask = 16'hBFFF;
defparam \addr_shift_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_shift_reg~9 (
	.dataa(\addr_shift_reg~7_combout ),
	.datab(\Equal1~0_combout ),
	.datac(sclk1),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\addr_shift_reg~9_combout ),
	.cout());
defparam \addr_shift_reg~9 .lut_mask = 16'hFFFE;
defparam \addr_shift_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_shift_reg~10 (
	.dataa(\next_addr[0]~q ),
	.datab(\addr_shift_reg~5_combout ),
	.datac(\Selector1~0_combout ),
	.datad(\addr_shift_reg~9_combout ),
	.cin(gnd),
	.combout(\addr_shift_reg~10_combout ),
	.cout());
defparam \addr_shift_reg~10 .lut_mask = 16'hFFFE;
defparam \addr_shift_reg~10 .sum_lutc_input = "datac";

dffeas \addr_shift_reg[0] (
	.clk(clock),
	.d(\addr_shift_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\addr_shift_reg[0]~q ),
	.prn(vcc));
defparam \addr_shift_reg[0] .is_wysiwyg = "true";
defparam \addr_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \addr_shift_reg~7 (
	.dataa(\addr_shift_reg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\currState.pauseState~q ),
	.cin(gnd),
	.combout(\addr_shift_reg~7_combout ),
	.cout());
defparam \addr_shift_reg~7 .lut_mask = 16'hAAFF;
defparam \addr_shift_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_shift_reg~8 (
	.dataa(\addr_shift_reg~7_combout ),
	.datab(\next_addr[1]~q ),
	.datac(\addr_shift_reg~5_combout ),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\addr_shift_reg~8_combout ),
	.cout());
defparam \addr_shift_reg~8 .lut_mask = 16'hFEFF;
defparam \addr_shift_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_shift_reg[3]~1 (
	.dataa(sclk1),
	.datab(\Equal1~3_combout ),
	.datac(\currState.pauseState~q ),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\addr_shift_reg[3]~1_combout ),
	.cout());
defparam \addr_shift_reg[3]~1 .lut_mask = 16'hFFF7;
defparam \addr_shift_reg[3]~1 .sum_lutc_input = "datac";

dffeas \addr_shift_reg[1] (
	.clk(clock),
	.d(\addr_shift_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\addr_shift_reg[3]~1_combout ),
	.q(\addr_shift_reg[1]~q ),
	.prn(vcc));
defparam \addr_shift_reg[1] .is_wysiwyg = "true";
defparam \addr_shift_reg[1] .power_up = "low";

cycloneive_lcell_comb \addr_shift_reg~4 (
	.dataa(\addr_shift_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\currState.pauseState~q ),
	.cin(gnd),
	.combout(\addr_shift_reg~4_combout ),
	.cout());
defparam \addr_shift_reg~4 .lut_mask = 16'hAAFF;
defparam \addr_shift_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_shift_reg~6 (
	.dataa(\addr_shift_reg~4_combout ),
	.datab(\next_addr[2]~q ),
	.datac(\addr_shift_reg~5_combout ),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\addr_shift_reg~6_combout ),
	.cout());
defparam \addr_shift_reg~6 .lut_mask = 16'hFEFF;
defparam \addr_shift_reg~6 .sum_lutc_input = "datac";

dffeas \addr_shift_reg[2] (
	.clk(clock),
	.d(\addr_shift_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\addr_shift_reg[3]~1_combout ),
	.q(\addr_shift_reg[2]~q ),
	.prn(vcc));
defparam \addr_shift_reg[2] .is_wysiwyg = "true";
defparam \addr_shift_reg[2] .power_up = "low";

cycloneive_lcell_comb \addr_shift_reg~3 (
	.dataa(\addr_shift_reg[2]~q ),
	.datab(go),
	.datac(\currState.waitState~q ),
	.datad(\currState.pauseState~q ),
	.cin(gnd),
	.combout(\addr_shift_reg~3_combout ),
	.cout());
defparam \addr_shift_reg~3 .lut_mask = 16'hBFFF;
defparam \addr_shift_reg~3 .sum_lutc_input = "datac";

dffeas \addr_shift_reg[3] (
	.clk(clock),
	.d(\addr_shift_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\addr_shift_reg[3]~1_combout ),
	.q(\addr_shift_reg[3]~q ),
	.prn(vcc));
defparam \addr_shift_reg[3] .is_wysiwyg = "true";
defparam \addr_shift_reg[3] .power_up = "low";

cycloneive_lcell_comb \addr_shift_reg~2 (
	.dataa(\addr_shift_reg[3]~q ),
	.datab(go),
	.datac(\currState.waitState~q ),
	.datad(\currState.pauseState~q ),
	.cin(gnd),
	.combout(\addr_shift_reg~2_combout ),
	.cout());
defparam \addr_shift_reg~2 .lut_mask = 16'hBFFF;
defparam \addr_shift_reg~2 .sum_lutc_input = "datac";

dffeas \addr_shift_reg[4] (
	.clk(clock),
	.d(\addr_shift_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\addr_shift_reg[3]~1_combout ),
	.q(\addr_shift_reg[4]~q ),
	.prn(vcc));
defparam \addr_shift_reg[4] .is_wysiwyg = "true";
defparam \addr_shift_reg[4] .power_up = "low";

cycloneive_lcell_comb \addr_shift_reg~0 (
	.dataa(\addr_shift_reg[4]~q ),
	.datab(go),
	.datac(\currState.waitState~q ),
	.datad(\currState.pauseState~q ),
	.cin(gnd),
	.combout(\addr_shift_reg~0_combout ),
	.cout());
defparam \addr_shift_reg~0 .lut_mask = 16'hBFFF;
defparam \addr_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\currState.pauseState~q ),
	.datab(\address[2]~q ),
	.datac(\address[1]~q ),
	.datad(\address[0]~q ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hBFFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~1 (
	.dataa(\Selector2~0_combout ),
	.datab(go),
	.datac(currStatedoneState),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
defparam \Selector2~1 .lut_mask = 16'hFEFE;
defparam \Selector2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~12 (
	.dataa(\address[1]~q ),
	.datab(\address[0]~q ),
	.datac(sclk1),
	.datad(\sclk_counter[3]~q ),
	.cin(gnd),
	.combout(\Decoder0~12_combout ),
	.cout());
defparam \Decoder0~12 .lut_mask = 16'hFFFE;
defparam \Decoder0~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~2 (
	.dataa(\address[2]~q ),
	.datab(\always5~0_combout ),
	.datac(\Equal1~3_combout ),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
defparam \Decoder0~2 .lut_mask = 16'hFFEF;
defparam \Decoder0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~3 (
	.dataa(\address[0]~q ),
	.datab(sclk1),
	.datac(\sclk_counter[3]~q ),
	.datad(\always5~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~3_combout ),
	.cout());
defparam \Decoder0~3 .lut_mask = 16'hFFFD;
defparam \Decoder0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~4 (
	.dataa(\address[2]~q ),
	.datab(\address[1]~q ),
	.datac(\Equal1~3_combout ),
	.datad(\Decoder0~3_combout ),
	.cin(gnd),
	.combout(\Decoder0~4_combout ),
	.cout());
defparam \Decoder0~4 .lut_mask = 16'hFFEF;
defparam \Decoder0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~5 (
	.dataa(\address[1]~q ),
	.datab(sclk1),
	.datac(\sclk_counter[3]~q ),
	.datad(\always5~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~5_combout ),
	.cout());
defparam \Decoder0~5 .lut_mask = 16'hFFFD;
defparam \Decoder0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~6 (
	.dataa(\address[2]~q ),
	.datab(\address[0]~q ),
	.datac(\Equal1~3_combout ),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~6_combout ),
	.cout());
defparam \Decoder0~6 .lut_mask = 16'hFFEF;
defparam \Decoder0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \reading7[6]~0 (
	.dataa(\address[2]~q ),
	.datab(\address[1]~q ),
	.datac(\Equal1~3_combout ),
	.datad(\Decoder0~3_combout ),
	.cin(gnd),
	.combout(\reading7[6]~0_combout ),
	.cout());
defparam \reading7[6]~0 .lut_mask = 16'hFF7F;
defparam \reading7[6]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~7 (
	.dataa(\address[2]~q ),
	.datab(sclk1),
	.datac(\sclk_counter[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~7_combout ),
	.cout());
defparam \Decoder0~7 .lut_mask = 16'hFDFD;
defparam \Decoder0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~8 (
	.dataa(\Add5~0_combout ),
	.datab(\always5~0_combout ),
	.datac(\Equal1~3_combout ),
	.datad(\Decoder0~7_combout ),
	.cin(gnd),
	.combout(\Decoder0~8_combout ),
	.cout());
defparam \Decoder0~8 .lut_mask = 16'hFFEF;
defparam \Decoder0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~9 (
	.dataa(\address[1]~q ),
	.datab(\address[2]~q ),
	.datac(\Equal1~3_combout ),
	.datad(\Decoder0~3_combout ),
	.cin(gnd),
	.combout(\Decoder0~9_combout ),
	.cout());
defparam \Decoder0~9 .lut_mask = 16'hFFBF;
defparam \Decoder0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~10 (
	.dataa(\address[0]~q ),
	.datab(\address[2]~q ),
	.datac(\Equal1~3_combout ),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~10_combout ),
	.cout());
defparam \Decoder0~10 .lut_mask = 16'hFFBF;
defparam \Decoder0~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~11 (
	.dataa(\always5~1_combout ),
	.datab(\address[2]~q ),
	.datac(\address[1]~q ),
	.datad(\address[0]~q ),
	.cin(gnd),
	.combout(\Decoder0~11_combout ),
	.cout());
defparam \Decoder0~11 .lut_mask = 16'hEFFF;
defparam \Decoder0~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always7~0 (
	.dataa(\Equal1~3_combout ),
	.datab(\sclk_counter[3]~q ),
	.datac(\always5~0_combout ),
	.datad(sclk1),
	.cin(gnd),
	.combout(\always7~0_combout ),
	.cout());
defparam \always7~0 .lut_mask = 16'hFF7F;
defparam \always7~0 .sum_lutc_input = "datac";

dffeas \shift_reg[0] (
	.clk(clock),
	.d(dout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[0]~q ),
	.prn(vcc));
defparam \shift_reg[0] .is_wysiwyg = "true";
defparam \shift_reg[0] .power_up = "low";

dffeas \shift_reg[1] (
	.clk(clock),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[1]~q ),
	.prn(vcc));
defparam \shift_reg[1] .is_wysiwyg = "true";
defparam \shift_reg[1] .power_up = "low";

dffeas \shift_reg[2] (
	.clk(clock),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[2]~q ),
	.prn(vcc));
defparam \shift_reg[2] .is_wysiwyg = "true";
defparam \shift_reg[2] .power_up = "low";

dffeas \shift_reg[3] (
	.clk(clock),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[3]~q ),
	.prn(vcc));
defparam \shift_reg[3] .is_wysiwyg = "true";
defparam \shift_reg[3] .power_up = "low";

dffeas \shift_reg[4] (
	.clk(clock),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[4]~q ),
	.prn(vcc));
defparam \shift_reg[4] .is_wysiwyg = "true";
defparam \shift_reg[4] .power_up = "low";

dffeas \shift_reg[5] (
	.clk(clock),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[5]~q ),
	.prn(vcc));
defparam \shift_reg[5] .is_wysiwyg = "true";
defparam \shift_reg[5] .power_up = "low";

dffeas \shift_reg[6] (
	.clk(clock),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[6]~q ),
	.prn(vcc));
defparam \shift_reg[6] .is_wysiwyg = "true";
defparam \shift_reg[6] .power_up = "low";

dffeas \shift_reg[7] (
	.clk(clock),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[7]~q ),
	.prn(vcc));
defparam \shift_reg[7] .is_wysiwyg = "true";
defparam \shift_reg[7] .power_up = "low";

dffeas \shift_reg[8] (
	.clk(clock),
	.d(\shift_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[8]~q ),
	.prn(vcc));
defparam \shift_reg[8] .is_wysiwyg = "true";
defparam \shift_reg[8] .power_up = "low";

dffeas \shift_reg[9] (
	.clk(clock),
	.d(\shift_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[9]~q ),
	.prn(vcc));
defparam \shift_reg[9] .is_wysiwyg = "true";
defparam \shift_reg[9] .power_up = "low";

dffeas \shift_reg[10] (
	.clk(clock),
	.d(\shift_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\shift_reg[10]~q ),
	.prn(vcc));
defparam \shift_reg[10] .is_wysiwyg = "true";
defparam \shift_reg[10] .power_up = "low";

endmodule

module niosII_niosII_cpu (
	wire_pll7_clk_0,
	sr_0,
	W_alu_result_6,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_5,
	W_alu_result_7,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	irq,
	irq1,
	readdata_4,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	d_read,
	d_write,
	d_writedata_0,
	d_byteenable_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_byteenable_1,
	i_read,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_8,
	F_pc_9,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	mem_84_0,
	mem_66_0,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	mem_54_0,
	src0_valid,
	WideOr1,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	d_writedata_10,
	d_byteenable_2,
	d_byteenable_3,
	src1_valid,
	read_accepted,
	src1_valid1,
	hbreak_enabled,
	d_writedata_8,
	d_writedata_9,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	WideOr11,
	rf_source_valid,
	uav_write,
	out_valid,
	av_readdata_pre_0,
	out_data_buffer_0,
	data_reg_0,
	out_payload_0,
	source_addr_1,
	F_iw_0,
	av_readdata_pre_1,
	out_data_buffer_1,
	out_payload_1,
	src_data_1,
	av_readdata_pre_2,
	out_data_buffer_2,
	data_reg_2,
	out_payload_2,
	F_iw_2,
	av_readdata_pre_3,
	out_data_buffer_3,
	out_payload_3,
	src_data_3,
	av_readdata_pre_4,
	out_data_buffer_4,
	out_payload_4,
	src_data_4,
	r_early_rst,
	src_data_46,
	av_readdata_pre_11,
	out_data_buffer_11,
	out_payload_11,
	src_data_11,
	av_readdata_pre_13,
	out_data_buffer_13,
	out_payload_13,
	src_data_13,
	av_readdata_pre_16,
	out_data_buffer_16,
	src_payload,
	av_readdata_pre_12,
	out_data_buffer_12,
	data_reg_12,
	out_payload_12,
	F_iw_12,
	av_readdata_pre_5,
	out_data_buffer_5,
	out_payload_5,
	src_data_5,
	av_readdata_pre_14,
	out_data_buffer_14,
	data_reg_14,
	out_payload_14,
	F_iw_14,
	av_readdata_pre_15,
	out_data_buffer_15,
	out_payload_15,
	src_data_15,
	av_readdata_pre_10,
	out_data_buffer_10,
	data_reg_10,
	out_payload_10,
	F_iw_10,
	av_readdata_pre_9,
	out_data_buffer_9,
	data_reg_9,
	out_payload_9,
	F_iw_9,
	av_readdata_pre_8,
	out_data_buffer_8,
	data_reg_8,
	out_payload_8,
	F_iw_8,
	av_readdata_pre_7,
	out_data_buffer_7,
	data_reg_7,
	out_payload_7,
	F_iw_7,
	av_readdata_pre_6,
	out_data_buffer_6,
	data_reg_6,
	out_payload_6,
	F_iw_6,
	av_readdata_pre_21,
	out_data_buffer_21,
	av_readdata_pre_30,
	out_data_buffer_30,
	av_readdata_pre_29,
	out_data_buffer_29,
	av_readdata_pre_28,
	out_data_buffer_28,
	av_readdata_pre_27,
	out_data_buffer_27,
	av_readdata_pre_26,
	out_data_buffer_26,
	av_readdata_pre_25,
	out_data_buffer_25,
	av_readdata_pre_24,
	out_data_buffer_24,
	av_readdata_pre_23,
	out_data_buffer_23,
	av_readdata_pre_22,
	out_data_buffer_22,
	av_readdata_pre_20,
	out_data_buffer_20,
	av_readdata_pre_19,
	out_data_buffer_19,
	av_readdata_pre_18,
	out_data_buffer_18,
	av_readdata_pre_17,
	out_data_buffer_17,
	out_valid1,
	src_data_0,
	dreg_1,
	timeout_occurred,
	control_register_0,
	dreg_11,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	src_data_12,
	src_data_2,
	src_data_21,
	src_data_31,
	av_readdata_pre_301,
	src_data_41,
	src_data_51,
	src_data_6,
	src_data_7,
	src_payload1,
	src_payload2,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_411,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_14,
	readdata_15,
	readdata_10,
	av_readdata_pre_31,
	out_data_buffer_31,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_6,
	readdata_26,
	out_data_buffer_261,
	readdata_21,
	readdata_30,
	readdata_25,
	out_data_buffer_251,
	src_payload3,
	readdata_29,
	readdata_24,
	out_data_buffer_241,
	readdata_28,
	src_payload4,
	readdata_27,
	src_payload5,
	readdata_261,
	src_payload6,
	readdata_251,
	src_payload7,
	readdata_241,
	src_payload8,
	readdata_23,
	src_payload9,
	readdata_22,
	src_payload10,
	src_payload11,
	readdata_20,
	src_data_151,
	readdata_19,
	src_data_14,
	readdata_18,
	src_data_131,
	readdata_17,
	src_data_121,
	src_data_111,
	src_data_10,
	src_data_9,
	src_data_8,
	src_payload12,
	readdata_271,
	out_data_buffer_271,
	readdata_281,
	out_data_buffer_281,
	readdata_291,
	out_data_buffer_291,
	readdata_301,
	out_data_buffer_301,
	readdata_31,
	out_data_buffer_311,
	readdata_311,
	debug_reset_request,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_data_33,
	src_payload17,
	src_payload18,
	src_data_34,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_data_35,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	sr_0;
output 	W_alu_result_6;
output 	W_alu_result_26;
output 	W_alu_result_25;
output 	W_alu_result_24;
output 	W_alu_result_23;
output 	W_alu_result_22;
output 	W_alu_result_21;
output 	W_alu_result_20;
output 	W_alu_result_19;
output 	W_alu_result_18;
output 	W_alu_result_17;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_12;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_5;
output 	W_alu_result_7;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_4;
output 	W_alu_result_3;
output 	W_alu_result_2;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
input 	irq;
input 	irq1;
output 	readdata_4;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
output 	d_read;
output 	d_write;
output 	d_writedata_0;
output 	d_byteenable_0;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
output 	d_byteenable_1;
output 	i_read;
output 	F_pc_24;
output 	F_pc_23;
output 	F_pc_22;
output 	F_pc_21;
output 	F_pc_20;
output 	F_pc_19;
output 	F_pc_18;
output 	F_pc_17;
output 	F_pc_16;
output 	F_pc_15;
output 	F_pc_14;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	F_pc_10;
output 	F_pc_8;
output 	F_pc_9;
output 	F_pc_0;
output 	F_pc_1;
output 	F_pc_2;
output 	F_pc_3;
output 	F_pc_4;
output 	F_pc_5;
output 	F_pc_6;
output 	F_pc_7;
input 	mem_84_0;
input 	mem_66_0;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	mem_54_0;
input 	src0_valid;
input 	WideOr1;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
output 	d_writedata_10;
output 	d_byteenable_2;
output 	d_byteenable_3;
input 	src1_valid;
input 	read_accepted;
input 	src1_valid1;
output 	hbreak_enabled;
output 	d_writedata_8;
output 	d_writedata_9;
output 	d_writedata_11;
output 	d_writedata_12;
output 	d_writedata_13;
output 	d_writedata_14;
output 	d_writedata_15;
output 	d_writedata_16;
output 	d_writedata_17;
output 	d_writedata_18;
output 	d_writedata_19;
output 	d_writedata_20;
output 	d_writedata_21;
output 	d_writedata_22;
output 	d_writedata_23;
input 	WideOr11;
input 	rf_source_valid;
input 	uav_write;
input 	out_valid;
input 	av_readdata_pre_0;
input 	out_data_buffer_0;
input 	data_reg_0;
input 	out_payload_0;
input 	source_addr_1;
output 	F_iw_0;
input 	av_readdata_pre_1;
input 	out_data_buffer_1;
input 	out_payload_1;
input 	src_data_1;
input 	av_readdata_pre_2;
input 	out_data_buffer_2;
input 	data_reg_2;
input 	out_payload_2;
output 	F_iw_2;
input 	av_readdata_pre_3;
input 	out_data_buffer_3;
input 	out_payload_3;
input 	src_data_3;
input 	av_readdata_pre_4;
input 	out_data_buffer_4;
input 	out_payload_4;
input 	src_data_4;
input 	r_early_rst;
input 	src_data_46;
input 	av_readdata_pre_11;
input 	out_data_buffer_11;
input 	out_payload_11;
input 	src_data_11;
input 	av_readdata_pre_13;
input 	out_data_buffer_13;
input 	out_payload_13;
input 	src_data_13;
input 	av_readdata_pre_16;
input 	out_data_buffer_16;
input 	src_payload;
input 	av_readdata_pre_12;
input 	out_data_buffer_12;
input 	data_reg_12;
input 	out_payload_12;
output 	F_iw_12;
input 	av_readdata_pre_5;
input 	out_data_buffer_5;
input 	out_payload_5;
input 	src_data_5;
input 	av_readdata_pre_14;
input 	out_data_buffer_14;
input 	data_reg_14;
input 	out_payload_14;
output 	F_iw_14;
input 	av_readdata_pre_15;
input 	out_data_buffer_15;
input 	out_payload_15;
input 	src_data_15;
input 	av_readdata_pre_10;
input 	out_data_buffer_10;
input 	data_reg_10;
input 	out_payload_10;
output 	F_iw_10;
input 	av_readdata_pre_9;
input 	out_data_buffer_9;
input 	data_reg_9;
input 	out_payload_9;
output 	F_iw_9;
input 	av_readdata_pre_8;
input 	out_data_buffer_8;
input 	data_reg_8;
input 	out_payload_8;
output 	F_iw_8;
input 	av_readdata_pre_7;
input 	out_data_buffer_7;
input 	data_reg_7;
input 	out_payload_7;
output 	F_iw_7;
input 	av_readdata_pre_6;
input 	out_data_buffer_6;
input 	data_reg_6;
input 	out_payload_6;
output 	F_iw_6;
input 	av_readdata_pre_21;
input 	out_data_buffer_21;
input 	av_readdata_pre_30;
input 	out_data_buffer_30;
input 	av_readdata_pre_29;
input 	out_data_buffer_29;
input 	av_readdata_pre_28;
input 	out_data_buffer_28;
input 	av_readdata_pre_27;
input 	out_data_buffer_27;
input 	av_readdata_pre_26;
input 	out_data_buffer_26;
input 	av_readdata_pre_25;
input 	out_data_buffer_25;
input 	av_readdata_pre_24;
input 	out_data_buffer_24;
input 	av_readdata_pre_23;
input 	out_data_buffer_23;
input 	av_readdata_pre_22;
input 	out_data_buffer_22;
input 	av_readdata_pre_20;
input 	out_data_buffer_20;
input 	av_readdata_pre_19;
input 	out_data_buffer_19;
input 	av_readdata_pre_18;
input 	out_data_buffer_18;
input 	av_readdata_pre_17;
input 	out_data_buffer_17;
input 	out_valid1;
input 	src_data_0;
input 	dreg_1;
input 	timeout_occurred;
input 	control_register_0;
input 	dreg_11;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
input 	src_data_12;
input 	src_data_2;
input 	src_data_21;
input 	src_data_31;
input 	av_readdata_pre_301;
input 	src_data_41;
input 	src_data_51;
input 	src_data_6;
input 	src_data_7;
input 	src_payload1;
input 	src_payload2;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_411;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_5;
output 	readdata_14;
output 	readdata_15;
output 	readdata_10;
input 	av_readdata_pre_31;
input 	out_data_buffer_31;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_6;
input 	readdata_26;
input 	out_data_buffer_261;
output 	readdata_21;
output 	readdata_30;
input 	readdata_25;
input 	out_data_buffer_251;
input 	src_payload3;
output 	readdata_29;
input 	readdata_24;
input 	out_data_buffer_241;
output 	readdata_28;
input 	src_payload4;
output 	readdata_27;
input 	src_payload5;
output 	readdata_261;
input 	src_payload6;
output 	readdata_251;
input 	src_payload7;
output 	readdata_241;
input 	src_payload8;
output 	readdata_23;
input 	src_payload9;
output 	readdata_22;
input 	src_payload10;
input 	src_payload11;
output 	readdata_20;
input 	src_data_151;
output 	readdata_19;
input 	src_data_14;
output 	readdata_18;
input 	src_data_131;
output 	readdata_17;
input 	src_data_121;
input 	src_data_111;
input 	src_data_10;
input 	src_data_9;
input 	src_data_8;
input 	src_payload12;
input 	readdata_271;
input 	out_data_buffer_271;
input 	readdata_281;
input 	out_data_buffer_281;
input 	readdata_291;
input 	out_data_buffer_291;
input 	readdata_301;
input 	out_data_buffer_301;
input 	readdata_31;
input 	out_data_buffer_311;
output 	readdata_311;
output 	debug_reset_request;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_data_33;
input 	src_payload17;
input 	src_payload18;
input 	src_data_34;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_data_35;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_niosII_cpu_cpu cpu(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.sr_0(sr_0),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.irq(irq),
	.irq1(irq1),
	.readdata_4(readdata_4),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.r_sync_rst(r_sync_rst),
	.d_read1(d_read),
	.d_write1(d_write),
	.d_writedata_0(d_writedata_0),
	.d_byteenable_0(d_byteenable_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_byteenable_1(d_byteenable_1),
	.i_read1(i_read),
	.F_pc_24(F_pc_24),
	.F_pc_23(F_pc_23),
	.F_pc_22(F_pc_22),
	.F_pc_21(F_pc_21),
	.F_pc_20(F_pc_20),
	.F_pc_19(F_pc_19),
	.F_pc_18(F_pc_18),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.F_pc_10(F_pc_10),
	.F_pc_8(F_pc_8),
	.F_pc_9(F_pc_9),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_7(F_pc_7),
	.mem_84_0(mem_84_0),
	.mem_66_0(mem_66_0),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.read_latency_shift_reg_02(read_latency_shift_reg_02),
	.mem_54_0(mem_54_0),
	.src0_valid(src0_valid),
	.WideOr1(WideOr1),
	.saved_grant_0(saved_grant_0),
	.debug_mem_slave_waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.av_waitrequest(av_waitrequest),
	.d_writedata_10(d_writedata_10),
	.d_byteenable_2(d_byteenable_2),
	.d_byteenable_3(d_byteenable_3),
	.src1_valid(src1_valid),
	.read_accepted(read_accepted),
	.src1_valid1(src1_valid1),
	.hbreak_enabled1(hbreak_enabled),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.WideOr11(WideOr11),
	.rf_source_valid(rf_source_valid),
	.uav_write(uav_write),
	.out_valid(out_valid),
	.av_readdata_pre_0(av_readdata_pre_0),
	.out_data_buffer_0(out_data_buffer_0),
	.data_reg_0(data_reg_0),
	.out_payload_0(out_payload_0),
	.source_addr_1(source_addr_1),
	.F_iw_0(F_iw_0),
	.av_readdata_pre_1(av_readdata_pre_1),
	.out_data_buffer_1(out_data_buffer_1),
	.out_payload_1(out_payload_1),
	.src_data_1(src_data_1),
	.av_readdata_pre_2(av_readdata_pre_2),
	.out_data_buffer_2(out_data_buffer_2),
	.data_reg_2(data_reg_2),
	.out_payload_2(out_payload_2),
	.F_iw_2(F_iw_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.out_data_buffer_3(out_data_buffer_3),
	.out_payload_3(out_payload_3),
	.src_data_3(src_data_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.out_data_buffer_4(out_data_buffer_4),
	.out_payload_4(out_payload_4),
	.src_data_4(src_data_4),
	.r_early_rst(r_early_rst),
	.src_data_46(src_data_46),
	.av_readdata_pre_11(av_readdata_pre_11),
	.out_data_buffer_11(out_data_buffer_11),
	.out_payload_11(out_payload_11),
	.src_data_11(src_data_11),
	.av_readdata_pre_13(av_readdata_pre_13),
	.out_data_buffer_13(out_data_buffer_13),
	.out_payload_13(out_payload_13),
	.src_data_13(src_data_13),
	.av_readdata_pre_16(av_readdata_pre_16),
	.out_data_buffer_16(out_data_buffer_16),
	.src_payload(src_payload),
	.av_readdata_pre_12(av_readdata_pre_12),
	.out_data_buffer_12(out_data_buffer_12),
	.data_reg_12(data_reg_12),
	.out_payload_12(out_payload_12),
	.F_iw_12(F_iw_12),
	.av_readdata_pre_5(av_readdata_pre_5),
	.out_data_buffer_5(out_data_buffer_5),
	.out_payload_5(out_payload_5),
	.src_data_5(src_data_5),
	.av_readdata_pre_14(av_readdata_pre_14),
	.out_data_buffer_14(out_data_buffer_14),
	.data_reg_14(data_reg_14),
	.out_payload_14(out_payload_14),
	.F_iw_14(F_iw_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.out_data_buffer_15(out_data_buffer_15),
	.out_payload_15(out_payload_15),
	.src_data_15(src_data_15),
	.av_readdata_pre_10(av_readdata_pre_10),
	.out_data_buffer_10(out_data_buffer_10),
	.data_reg_10(data_reg_10),
	.out_payload_10(out_payload_10),
	.F_iw_10(F_iw_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.out_data_buffer_9(out_data_buffer_9),
	.data_reg_9(data_reg_9),
	.out_payload_9(out_payload_9),
	.F_iw_9(F_iw_9),
	.av_readdata_pre_8(av_readdata_pre_8),
	.out_data_buffer_8(out_data_buffer_8),
	.data_reg_8(data_reg_8),
	.out_payload_8(out_payload_8),
	.F_iw_8(F_iw_8),
	.av_readdata_pre_7(av_readdata_pre_7),
	.out_data_buffer_7(out_data_buffer_7),
	.data_reg_7(data_reg_7),
	.out_payload_7(out_payload_7),
	.F_iw_7(F_iw_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.out_data_buffer_6(out_data_buffer_6),
	.data_reg_6(data_reg_6),
	.out_payload_6(out_payload_6),
	.F_iw_6(F_iw_6),
	.av_readdata_pre_21(av_readdata_pre_21),
	.out_data_buffer_21(out_data_buffer_21),
	.av_readdata_pre_30(av_readdata_pre_30),
	.out_data_buffer_30(out_data_buffer_30),
	.av_readdata_pre_29(av_readdata_pre_29),
	.out_data_buffer_29(out_data_buffer_29),
	.av_readdata_pre_28(av_readdata_pre_28),
	.out_data_buffer_28(out_data_buffer_28),
	.av_readdata_pre_27(av_readdata_pre_27),
	.out_data_buffer_27(out_data_buffer_27),
	.av_readdata_pre_26(av_readdata_pre_26),
	.out_data_buffer_26(out_data_buffer_26),
	.av_readdata_pre_25(av_readdata_pre_25),
	.out_data_buffer_25(out_data_buffer_25),
	.av_readdata_pre_24(av_readdata_pre_24),
	.out_data_buffer_24(out_data_buffer_24),
	.av_readdata_pre_23(av_readdata_pre_23),
	.out_data_buffer_23(out_data_buffer_23),
	.av_readdata_pre_22(av_readdata_pre_22),
	.out_data_buffer_22(out_data_buffer_22),
	.av_readdata_pre_20(av_readdata_pre_20),
	.out_data_buffer_20(out_data_buffer_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.out_data_buffer_19(out_data_buffer_19),
	.av_readdata_pre_18(av_readdata_pre_18),
	.out_data_buffer_18(out_data_buffer_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.out_data_buffer_17(out_data_buffer_17),
	.out_valid1(out_valid1),
	.src_data_0(src_data_0),
	.dreg_1(dreg_1),
	.timeout_occurred(timeout_occurred),
	.control_register_0(control_register_0),
	.dreg_11(dreg_11),
	.readdata_0(readdata_0),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.readdata_3(readdata_3),
	.src_data_12(src_data_12),
	.src_data_2(src_data_2),
	.src_data_21(src_data_21),
	.src_data_31(src_data_31),
	.av_readdata_pre_301(av_readdata_pre_301),
	.src_data_41(src_data_41),
	.src_data_51(src_data_51),
	.src_data_6(src_data_6),
	.src_data_7(src_data_7),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_411(src_data_411),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_32(src_data_32),
	.readdata_11(readdata_11),
	.readdata_13(readdata_13),
	.readdata_16(readdata_16),
	.readdata_12(readdata_12),
	.readdata_5(readdata_5),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_10(readdata_10),
	.av_readdata_pre_31(av_readdata_pre_31),
	.out_data_buffer_31(out_data_buffer_31),
	.readdata_9(readdata_9),
	.readdata_8(readdata_8),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.readdata_26(readdata_26),
	.out_data_buffer_261(out_data_buffer_261),
	.readdata_21(readdata_21),
	.readdata_30(readdata_30),
	.readdata_25(readdata_25),
	.out_data_buffer_251(out_data_buffer_251),
	.src_payload3(src_payload3),
	.readdata_29(readdata_29),
	.readdata_24(readdata_24),
	.out_data_buffer_241(out_data_buffer_241),
	.readdata_28(readdata_28),
	.src_payload4(src_payload4),
	.readdata_27(readdata_27),
	.src_payload5(src_payload5),
	.readdata_261(readdata_261),
	.src_payload6(src_payload6),
	.readdata_251(readdata_251),
	.src_payload7(src_payload7),
	.readdata_241(readdata_241),
	.src_payload8(src_payload8),
	.readdata_23(readdata_23),
	.src_payload9(src_payload9),
	.readdata_22(readdata_22),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.readdata_20(readdata_20),
	.src_data_151(src_data_151),
	.readdata_19(readdata_19),
	.src_data_14(src_data_14),
	.readdata_18(readdata_18),
	.src_data_131(src_data_131),
	.readdata_17(readdata_17),
	.src_data_121(src_data_121),
	.src_data_111(src_data_111),
	.src_data_10(src_data_10),
	.src_data_9(src_data_9),
	.src_data_8(src_data_8),
	.src_payload12(src_payload12),
	.readdata_271(readdata_271),
	.out_data_buffer_271(out_data_buffer_271),
	.readdata_281(readdata_281),
	.out_data_buffer_281(out_data_buffer_281),
	.readdata_291(readdata_291),
	.out_data_buffer_291(out_data_buffer_291),
	.readdata_301(readdata_301),
	.out_data_buffer_301(out_data_buffer_301),
	.readdata_31(readdata_31),
	.out_data_buffer_311(out_data_buffer_311),
	.readdata_311(readdata_311),
	.debug_reset_request(debug_reset_request),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_data_33(src_data_33),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_data_34(src_data_34),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_data_35(src_data_35),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.src_payload32(src_payload32),
	.src_payload33(src_payload33),
	.src_payload34(src_payload34),
	.src_payload35(src_payload35),
	.src_payload36(src_payload36),
	.src_payload37(src_payload37),
	.src_payload38(src_payload38),
	.src_payload39(src_payload39),
	.src_payload40(src_payload40),
	.src_payload41(src_payload41),
	.src_payload42(src_payload42),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

endmodule

module niosII_niosII_cpu_cpu (
	wire_pll7_clk_0,
	sr_0,
	W_alu_result_6,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_5,
	W_alu_result_7,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	irq,
	irq1,
	readdata_4,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	d_read1,
	d_write1,
	d_writedata_0,
	d_byteenable_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_byteenable_1,
	i_read1,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_8,
	F_pc_9,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	mem_84_0,
	mem_66_0,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	mem_54_0,
	src0_valid,
	WideOr1,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	d_writedata_10,
	d_byteenable_2,
	d_byteenable_3,
	src1_valid,
	read_accepted,
	src1_valid1,
	hbreak_enabled1,
	d_writedata_8,
	d_writedata_9,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	WideOr11,
	rf_source_valid,
	uav_write,
	out_valid,
	av_readdata_pre_0,
	out_data_buffer_0,
	data_reg_0,
	out_payload_0,
	source_addr_1,
	F_iw_0,
	av_readdata_pre_1,
	out_data_buffer_1,
	out_payload_1,
	src_data_1,
	av_readdata_pre_2,
	out_data_buffer_2,
	data_reg_2,
	out_payload_2,
	F_iw_2,
	av_readdata_pre_3,
	out_data_buffer_3,
	out_payload_3,
	src_data_3,
	av_readdata_pre_4,
	out_data_buffer_4,
	out_payload_4,
	src_data_4,
	r_early_rst,
	src_data_46,
	av_readdata_pre_11,
	out_data_buffer_11,
	out_payload_11,
	src_data_11,
	av_readdata_pre_13,
	out_data_buffer_13,
	out_payload_13,
	src_data_13,
	av_readdata_pre_16,
	out_data_buffer_16,
	src_payload,
	av_readdata_pre_12,
	out_data_buffer_12,
	data_reg_12,
	out_payload_12,
	F_iw_12,
	av_readdata_pre_5,
	out_data_buffer_5,
	out_payload_5,
	src_data_5,
	av_readdata_pre_14,
	out_data_buffer_14,
	data_reg_14,
	out_payload_14,
	F_iw_14,
	av_readdata_pre_15,
	out_data_buffer_15,
	out_payload_15,
	src_data_15,
	av_readdata_pre_10,
	out_data_buffer_10,
	data_reg_10,
	out_payload_10,
	F_iw_10,
	av_readdata_pre_9,
	out_data_buffer_9,
	data_reg_9,
	out_payload_9,
	F_iw_9,
	av_readdata_pre_8,
	out_data_buffer_8,
	data_reg_8,
	out_payload_8,
	F_iw_8,
	av_readdata_pre_7,
	out_data_buffer_7,
	data_reg_7,
	out_payload_7,
	F_iw_7,
	av_readdata_pre_6,
	out_data_buffer_6,
	data_reg_6,
	out_payload_6,
	F_iw_6,
	av_readdata_pre_21,
	out_data_buffer_21,
	av_readdata_pre_30,
	out_data_buffer_30,
	av_readdata_pre_29,
	out_data_buffer_29,
	av_readdata_pre_28,
	out_data_buffer_28,
	av_readdata_pre_27,
	out_data_buffer_27,
	av_readdata_pre_26,
	out_data_buffer_26,
	av_readdata_pre_25,
	out_data_buffer_25,
	av_readdata_pre_24,
	out_data_buffer_24,
	av_readdata_pre_23,
	out_data_buffer_23,
	av_readdata_pre_22,
	out_data_buffer_22,
	av_readdata_pre_20,
	out_data_buffer_20,
	av_readdata_pre_19,
	out_data_buffer_19,
	av_readdata_pre_18,
	out_data_buffer_18,
	av_readdata_pre_17,
	out_data_buffer_17,
	out_valid1,
	src_data_0,
	dreg_1,
	timeout_occurred,
	control_register_0,
	dreg_11,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	src_data_12,
	src_data_2,
	src_data_21,
	src_data_31,
	av_readdata_pre_301,
	src_data_41,
	src_data_51,
	src_data_6,
	src_data_7,
	src_payload1,
	src_payload2,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_411,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_14,
	readdata_15,
	readdata_10,
	av_readdata_pre_31,
	out_data_buffer_31,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_6,
	readdata_26,
	out_data_buffer_261,
	readdata_21,
	readdata_30,
	readdata_25,
	out_data_buffer_251,
	src_payload3,
	readdata_29,
	readdata_24,
	out_data_buffer_241,
	readdata_28,
	src_payload4,
	readdata_27,
	src_payload5,
	readdata_261,
	src_payload6,
	readdata_251,
	src_payload7,
	readdata_241,
	src_payload8,
	readdata_23,
	src_payload9,
	readdata_22,
	src_payload10,
	src_payload11,
	readdata_20,
	src_data_151,
	readdata_19,
	src_data_14,
	readdata_18,
	src_data_131,
	readdata_17,
	src_data_121,
	src_data_111,
	src_data_10,
	src_data_9,
	src_data_8,
	src_payload12,
	readdata_271,
	out_data_buffer_271,
	readdata_281,
	out_data_buffer_281,
	readdata_291,
	out_data_buffer_291,
	readdata_301,
	out_data_buffer_301,
	readdata_31,
	out_data_buffer_311,
	readdata_311,
	debug_reset_request,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_data_33,
	src_payload17,
	src_payload18,
	src_data_34,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_data_35,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	sr_0;
output 	W_alu_result_6;
output 	W_alu_result_26;
output 	W_alu_result_25;
output 	W_alu_result_24;
output 	W_alu_result_23;
output 	W_alu_result_22;
output 	W_alu_result_21;
output 	W_alu_result_20;
output 	W_alu_result_19;
output 	W_alu_result_18;
output 	W_alu_result_17;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_12;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_5;
output 	W_alu_result_7;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_4;
output 	W_alu_result_3;
output 	W_alu_result_2;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
input 	irq;
input 	irq1;
output 	readdata_4;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
output 	d_read1;
output 	d_write1;
output 	d_writedata_0;
output 	d_byteenable_0;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
output 	d_byteenable_1;
output 	i_read1;
output 	F_pc_24;
output 	F_pc_23;
output 	F_pc_22;
output 	F_pc_21;
output 	F_pc_20;
output 	F_pc_19;
output 	F_pc_18;
output 	F_pc_17;
output 	F_pc_16;
output 	F_pc_15;
output 	F_pc_14;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	F_pc_10;
output 	F_pc_8;
output 	F_pc_9;
output 	F_pc_0;
output 	F_pc_1;
output 	F_pc_2;
output 	F_pc_3;
output 	F_pc_4;
output 	F_pc_5;
output 	F_pc_6;
output 	F_pc_7;
input 	mem_84_0;
input 	mem_66_0;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	mem_54_0;
input 	src0_valid;
input 	WideOr1;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
output 	d_writedata_10;
output 	d_byteenable_2;
output 	d_byteenable_3;
input 	src1_valid;
input 	read_accepted;
input 	src1_valid1;
output 	hbreak_enabled1;
output 	d_writedata_8;
output 	d_writedata_9;
output 	d_writedata_11;
output 	d_writedata_12;
output 	d_writedata_13;
output 	d_writedata_14;
output 	d_writedata_15;
output 	d_writedata_16;
output 	d_writedata_17;
output 	d_writedata_18;
output 	d_writedata_19;
output 	d_writedata_20;
output 	d_writedata_21;
output 	d_writedata_22;
output 	d_writedata_23;
input 	WideOr11;
input 	rf_source_valid;
input 	uav_write;
input 	out_valid;
input 	av_readdata_pre_0;
input 	out_data_buffer_0;
input 	data_reg_0;
input 	out_payload_0;
input 	source_addr_1;
output 	F_iw_0;
input 	av_readdata_pre_1;
input 	out_data_buffer_1;
input 	out_payload_1;
input 	src_data_1;
input 	av_readdata_pre_2;
input 	out_data_buffer_2;
input 	data_reg_2;
input 	out_payload_2;
output 	F_iw_2;
input 	av_readdata_pre_3;
input 	out_data_buffer_3;
input 	out_payload_3;
input 	src_data_3;
input 	av_readdata_pre_4;
input 	out_data_buffer_4;
input 	out_payload_4;
input 	src_data_4;
input 	r_early_rst;
input 	src_data_46;
input 	av_readdata_pre_11;
input 	out_data_buffer_11;
input 	out_payload_11;
input 	src_data_11;
input 	av_readdata_pre_13;
input 	out_data_buffer_13;
input 	out_payload_13;
input 	src_data_13;
input 	av_readdata_pre_16;
input 	out_data_buffer_16;
input 	src_payload;
input 	av_readdata_pre_12;
input 	out_data_buffer_12;
input 	data_reg_12;
input 	out_payload_12;
output 	F_iw_12;
input 	av_readdata_pre_5;
input 	out_data_buffer_5;
input 	out_payload_5;
input 	src_data_5;
input 	av_readdata_pre_14;
input 	out_data_buffer_14;
input 	data_reg_14;
input 	out_payload_14;
output 	F_iw_14;
input 	av_readdata_pre_15;
input 	out_data_buffer_15;
input 	out_payload_15;
input 	src_data_15;
input 	av_readdata_pre_10;
input 	out_data_buffer_10;
input 	data_reg_10;
input 	out_payload_10;
output 	F_iw_10;
input 	av_readdata_pre_9;
input 	out_data_buffer_9;
input 	data_reg_9;
input 	out_payload_9;
output 	F_iw_9;
input 	av_readdata_pre_8;
input 	out_data_buffer_8;
input 	data_reg_8;
input 	out_payload_8;
output 	F_iw_8;
input 	av_readdata_pre_7;
input 	out_data_buffer_7;
input 	data_reg_7;
input 	out_payload_7;
output 	F_iw_7;
input 	av_readdata_pre_6;
input 	out_data_buffer_6;
input 	data_reg_6;
input 	out_payload_6;
output 	F_iw_6;
input 	av_readdata_pre_21;
input 	out_data_buffer_21;
input 	av_readdata_pre_30;
input 	out_data_buffer_30;
input 	av_readdata_pre_29;
input 	out_data_buffer_29;
input 	av_readdata_pre_28;
input 	out_data_buffer_28;
input 	av_readdata_pre_27;
input 	out_data_buffer_27;
input 	av_readdata_pre_26;
input 	out_data_buffer_26;
input 	av_readdata_pre_25;
input 	out_data_buffer_25;
input 	av_readdata_pre_24;
input 	out_data_buffer_24;
input 	av_readdata_pre_23;
input 	out_data_buffer_23;
input 	av_readdata_pre_22;
input 	out_data_buffer_22;
input 	av_readdata_pre_20;
input 	out_data_buffer_20;
input 	av_readdata_pre_19;
input 	out_data_buffer_19;
input 	av_readdata_pre_18;
input 	out_data_buffer_18;
input 	av_readdata_pre_17;
input 	out_data_buffer_17;
input 	out_valid1;
input 	src_data_0;
input 	dreg_1;
input 	timeout_occurred;
input 	control_register_0;
input 	dreg_11;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
input 	src_data_12;
input 	src_data_2;
input 	src_data_21;
input 	src_data_31;
input 	av_readdata_pre_301;
input 	src_data_41;
input 	src_data_51;
input 	src_data_6;
input 	src_data_7;
input 	src_payload1;
input 	src_payload2;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_411;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_5;
output 	readdata_14;
output 	readdata_15;
output 	readdata_10;
input 	av_readdata_pre_31;
input 	out_data_buffer_31;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_6;
input 	readdata_26;
input 	out_data_buffer_261;
output 	readdata_21;
output 	readdata_30;
input 	readdata_25;
input 	out_data_buffer_251;
input 	src_payload3;
output 	readdata_29;
input 	readdata_24;
input 	out_data_buffer_241;
output 	readdata_28;
input 	src_payload4;
output 	readdata_27;
input 	src_payload5;
output 	readdata_261;
input 	src_payload6;
output 	readdata_251;
input 	src_payload7;
output 	readdata_241;
input 	src_payload8;
output 	readdata_23;
input 	src_payload9;
output 	readdata_22;
input 	src_payload10;
input 	src_payload11;
output 	readdata_20;
input 	src_data_151;
output 	readdata_19;
input 	src_data_14;
output 	readdata_18;
input 	src_data_131;
output 	readdata_17;
input 	src_data_121;
input 	src_data_111;
input 	src_data_10;
input 	src_data_9;
input 	src_data_8;
input 	src_payload12;
input 	readdata_271;
input 	out_data_buffer_271;
input 	readdata_281;
input 	out_data_buffer_281;
input 	readdata_291;
input 	out_data_buffer_291;
input 	readdata_301;
input 	out_data_buffer_301;
input 	readdata_31;
input 	out_data_buffer_311;
output 	readdata_311;
output 	debug_reset_request;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_data_33;
input 	src_payload17;
input 	src_payload18;
input 	src_data_34;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_data_35;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \W_alu_result[0]~q ;
wire \the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_oci_debug|jtag_break~q ;
wire \W_alu_result[1]~q ;
wire \Add1~88_combout ;
wire \Add1~90_combout ;
wire \Add1~92_combout ;
wire \Add1~94_combout ;
wire \Add1~96_combout ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \av_ld_byte2_data[7]~q ;
wire \av_ld_byte2_data[6]~q ;
wire \av_ld_byte2_data[5]~q ;
wire \av_ld_byte2_data[4]~q ;
wire \av_ld_byte2_data[3]~q ;
wire \av_ld_byte2_data[2]~q ;
wire \av_ld_byte2_data[1]~q ;
wire \av_ld_byte2_data[0]~q ;
wire \av_ld_byte1_data[7]~q ;
wire \av_ld_byte1_data[6]~q ;
wire \av_ld_byte1_data[5]~q ;
wire \av_ld_byte1_data[4]~q ;
wire \av_ld_byte1_data[3]~q ;
wire \av_ld_byte1_data[2]~q ;
wire \av_ld_byte1_data[1]~q ;
wire \av_ld_byte1_data[0]~q ;
wire \W_alu_result[0]~25_combout ;
wire \W_alu_result[1]~26_combout ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \W_alu_result[27]~q ;
wire \W_alu_result[28]~q ;
wire \W_alu_result[29]~q ;
wire \W_alu_result[30]~q ;
wire \W_alu_result[31]~q ;
wire \av_ld_byte2_data[7]~0_combout ;
wire \av_ld_byte2_data[6]~1_combout ;
wire \av_ld_byte2_data[5]~2_combout ;
wire \av_ld_byte2_data[4]~3_combout ;
wire \av_ld_byte2_data[3]~4_combout ;
wire \av_ld_byte2_data[2]~5_combout ;
wire \av_ld_byte2_data[1]~6_combout ;
wire \av_ld_byte2_data[0]~7_combout ;
wire \av_ld_byte1_data[7]~0_combout ;
wire \av_ld_byte1_data[6]~1_combout ;
wire \av_ld_byte1_data[5]~2_combout ;
wire \av_ld_byte1_data[4]~3_combout ;
wire \av_ld_byte1_data[3]~4_combout ;
wire \av_ld_byte1_data[2]~5_combout ;
wire \av_ld_byte1_data[1]~6_combout ;
wire \av_ld_byte1_data[0]~7_combout ;
wire \W_alu_result[27]~27_combout ;
wire \W_alu_result[28]~28_combout ;
wire \W_alu_result[29]~29_combout ;
wire \W_alu_result[30]~30_combout ;
wire \W_alu_result[31]~31_combout ;
wire \D_ctrl_ld_signed~1_combout ;
wire \R_wr_dst_reg~q ;
wire \W_rf_wren~combout ;
wire \av_ld_byte0_data[0]~q ;
wire \W_rf_wr_data[0]~0_combout ;
wire \W_control_rd_data[0]~q ;
wire \W_rf_wr_data[0]~1_combout ;
wire \W_rf_wr_data[0]~2_combout ;
wire \R_dst_regnum[0]~q ;
wire \R_dst_regnum[1]~q ;
wire \R_dst_regnum[2]~q ;
wire \R_dst_regnum[3]~q ;
wire \R_dst_regnum[4]~q ;
wire \av_ld_byte0_data[1]~q ;
wire \W_control_rd_data[1]~q ;
wire \W_rf_wr_data[1]~3_combout ;
wire \W_rf_wr_data[1]~4_combout ;
wire \av_ld_byte0_data[2]~q ;
wire \W_control_rd_data[2]~q ;
wire \W_rf_wr_data[2]~5_combout ;
wire \W_rf_wr_data[2]~6_combout ;
wire \av_ld_byte0_data[3]~q ;
wire \W_control_rd_data[3]~q ;
wire \W_rf_wr_data[3]~7_combout ;
wire \W_rf_wr_data[3]~8_combout ;
wire \av_ld_byte0_data[4]~q ;
wire \W_control_rd_data[4]~q ;
wire \W_rf_wr_data[4]~9_combout ;
wire \W_rf_wr_data[4]~10_combout ;
wire \av_ld_byte0_data[5]~q ;
wire \W_rf_wr_data[5]~11_combout ;
wire \av_ld_byte0_data[6]~q ;
wire \W_rf_wr_data[6]~12_combout ;
wire \av_ld_byte0_data[7]~q ;
wire \W_rf_wr_data[7]~13_combout ;
wire \D_iw[31]~q ;
wire \av_ld_byte3_data[2]~q ;
wire \W_rf_wr_data[26]~14_combout ;
wire \av_ld_byte3_data[1]~q ;
wire \W_rf_wr_data[25]~15_combout ;
wire \av_ld_byte3_data[0]~q ;
wire \W_rf_wr_data[24]~16_combout ;
wire \W_rf_wr_data[23]~17_combout ;
wire \W_rf_wr_data[22]~18_combout ;
wire \W_rf_wr_data[21]~19_combout ;
wire \W_rf_wr_data[20]~20_combout ;
wire \W_rf_wr_data[19]~21_combout ;
wire \W_rf_wr_data[18]~22_combout ;
wire \W_rf_wr_data[17]~23_combout ;
wire \W_rf_wr_data[16]~24_combout ;
wire \W_rf_wr_data[15]~25_combout ;
wire \W_rf_wr_data[14]~26_combout ;
wire \W_rf_wr_data[13]~27_combout ;
wire \W_rf_wr_data[12]~28_combout ;
wire \W_rf_wr_data[11]~29_combout ;
wire \W_rf_wr_data[10]~30_combout ;
wire \W_rf_wr_data[9]~31_combout ;
wire \W_rf_wr_data[8]~32_combout ;
wire \D_wr_dst_reg~0_combout ;
wire \D_wr_dst_reg~1_combout ;
wire \D_dst_regnum[1]~0_combout ;
wire \D_ctrl_implicit_dst_eretaddr~3_combout ;
wire \D_ctrl_implicit_dst_eretaddr~4_combout ;
wire \D_ctrl_implicit_dst_eretaddr~5_combout ;
wire \D_ctrl_implicit_dst_eretaddr~6_combout ;
wire \D_dst_regnum[1]~1_combout ;
wire \D_dst_regnum[2]~2_combout ;
wire \D_dst_regnum[2]~3_combout ;
wire \D_dst_regnum[2]~4_combout ;
wire \D_dst_regnum[2]~5_combout ;
wire \D_dst_regnum[4]~6_combout ;
wire \D_dst_regnum[3]~7_combout ;
wire \Equal0~19_combout ;
wire \D_dst_regnum[0]~8_combout ;
wire \D_wr_dst_reg~2_combout ;
wire \av_ld_rshift8~0_combout ;
wire \av_ld_rshift8~1_combout ;
wire \av_ld_byte0_data[2]~0_combout ;
wire \E_control_rd_data[0]~0_combout ;
wire \E_control_rd_data[0]~1_combout ;
wire \E_control_rd_data[0]~2_combout ;
wire \E_control_rd_data[0]~3_combout ;
wire \the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[4]~q ;
wire \the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[3]~q ;
wire \the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[2]~q ;
wire \the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[1]~q ;
wire \the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[0]~q ;
wire \the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ;
wire \W_control_rd_data[1]~0_combout ;
wire \E_control_rd_data[1]~4_combout ;
wire \av_ld_byte0_data_nxt[2]~14_combout ;
wire \E_control_rd_data[2]~5_combout ;
wire \E_control_rd_data[3]~6_combout ;
wire \E_control_rd_data[4]~7_combout ;
wire \av_ld_byte3_data[3]~q ;
wire \W_rf_wr_data[27]~33_combout ;
wire \av_ld_byte3_data[4]~q ;
wire \W_rf_wr_data[28]~34_combout ;
wire \av_ld_byte3_data[5]~q ;
wire \W_rf_wr_data[29]~35_combout ;
wire \av_ld_byte3_data[6]~q ;
wire \W_rf_wr_data[30]~36_combout ;
wire \av_ld_byte3_data[7]~q ;
wire \W_rf_wr_data[31]~37_combout ;
wire \F_iw[31]~76_combout ;
wire \F_iw[31]~77_combout ;
wire \R_ctrl_ld_signed~q ;
wire \av_fill_bit~0_combout ;
wire \av_ld_byte3_data_nxt~0_combout ;
wire \av_ld_byte3_data_nxt~1_combout ;
wire \av_ld_byte3_data_nxt~2_combout ;
wire \av_ld_byte3_data_nxt~3_combout ;
wire \av_ld_byte3_data_nxt~4_combout ;
wire \av_ld_byte3_data_nxt~5_combout ;
wire \av_ld_byte3_data_nxt~6_combout ;
wire \av_ld_byte3_data_nxt~7_combout ;
wire \av_ld_byte3_data_nxt~8_combout ;
wire \av_ld_byte3_data_nxt~9_combout ;
wire \av_ld_byte3_data_nxt~10_combout ;
wire \av_ld_byte3_data_nxt~11_combout ;
wire \av_ld_byte3_data_nxt~12_combout ;
wire \av_ld_byte1_data_en~0_combout ;
wire \av_ld_byte3_data_nxt~13_combout ;
wire \av_ld_byte3_data_nxt~14_combout ;
wire \av_ld_byte3_data_nxt~15_combout ;
wire \av_ld_byte3_data_nxt~16_combout ;
wire \av_ld_byte3_data_nxt~17_combout ;
wire \av_ld_byte3_data_nxt~18_combout ;
wire \av_ld_byte3_data_nxt~19_combout ;
wire \av_ld_byte3_data_nxt~20_combout ;
wire \av_ld_byte3_data_nxt~21_combout ;
wire \av_ld_byte3_data_nxt~22_combout ;
wire \av_ld_byte3_data_nxt~23_combout ;
wire \av_ld_byte3_data_nxt~24_combout ;
wire \av_ld_byte3_data_nxt~25_combout ;
wire \av_ld_byte3_data_nxt~26_combout ;
wire \av_ld_byte3_data_nxt~27_combout ;
wire \av_ld_byte3_data_nxt~28_combout ;
wire \av_ld_byte3_data_nxt~29_combout ;
wire \av_ld_byte3_data_nxt~30_combout ;
wire \av_ld_byte3_data_nxt~31_combout ;
wire \av_ld_byte3_data_nxt~32_combout ;
wire \av_ld_byte3_data_nxt~33_combout ;
wire \av_ld_byte3_data_nxt~34_combout ;
wire \av_ld_byte3_data_nxt~35_combout ;
wire \av_ld_byte0_data_nxt[0]~15_combout ;
wire \av_ld_byte0_data_nxt[1]~16_combout ;
wire \av_ld_byte0_data_nxt[3]~17_combout ;
wire \av_ld_byte0_data_nxt[4]~18_combout ;
wire \av_ld_byte0_data_nxt[5]~19_combout ;
wire \av_ld_byte0_data_nxt[6]~20_combout ;
wire \av_ld_byte0_data_nxt[7]~21_combout ;
wire \F_valid~0_combout ;
wire \D_valid~q ;
wire \R_valid~q ;
wire \F_iw[11]~16_combout ;
wire \F_iw[8]~38_combout ;
wire \F_iw[8]~40_combout ;
wire \D_iw[8]~q ;
wire \F_iw[4]~14_combout ;
wire \F_iw[4]~15_combout ;
wire \D_iw[4]~q ;
wire \F_iw[5]~25_combout ;
wire \F_iw[5]~26_combout ;
wire \D_iw[5]~q ;
wire \F_iw[0]~4_combout ;
wire \F_iw[0]~6_combout ;
wire \D_iw[0]~q ;
wire \F_iw[1]~7_combout ;
wire \F_iw[1]~8_combout ;
wire \D_iw[1]~q ;
wire \F_iw[3]~12_combout ;
wire \F_iw[3]~13_combout ;
wire \D_iw[3]~q ;
wire \F_iw[2]~9_combout ;
wire \F_iw[2]~11_combout ;
wire \D_iw[2]~q ;
wire \Equal0~7_combout ;
wire \Equal0~8_combout ;
wire \F_iw[15]~30_combout ;
wire \F_iw[15]~31_combout ;
wire \D_iw[15]~q ;
wire \E_new_inst~q ;
wire \D_ctrl_st~0_combout ;
wire \R_ctrl_st~q ;
wire \W_valid~3_combout ;
wire \W_valid~2_combout ;
wire \W_valid~q ;
wire \hbreak_pending_nxt~0_combout ;
wire \hbreak_pending~q ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \F_iw[14]~27_combout ;
wire \F_iw[14]~29_combout ;
wire \F_iw[14]~78_combout ;
wire \D_iw[14]~q ;
wire \D_op_opx_rsv63~0_combout ;
wire \F_iw[13]~18_combout ;
wire \F_iw[13]~19_combout ;
wire \D_iw[13]~q ;
wire \F_iw[16]~20_combout ;
wire \F_iw[16]~21_combout ;
wire \D_iw[16]~q ;
wire \F_iw[12]~22_combout ;
wire \F_iw[12]~24_combout ;
wire \D_iw[12]~q ;
wire \Equal62~4_combout ;
wire \Equal62~5_combout ;
wire \Equal62~6_combout ;
wire \D_ctrl_shift_rot~0_combout ;
wire \Equal62~7_combout ;
wire \D_ctrl_shift_rot~1_combout ;
wire \D_ctrl_shift_logical~0_combout ;
wire \D_ctrl_shift_rot~2_combout ;
wire \D_ctrl_shift_rot~3_combout ;
wire \R_ctrl_shift_rot~q ;
wire \E_shift_rot_cnt[0]~5_combout ;
wire \D_ctrl_hi_imm16~0_combout ;
wire \D_ctrl_hi_imm16~1_combout ;
wire \R_ctrl_hi_imm16~q ;
wire \Equal0~14_combout ;
wire \D_ctrl_alu_force_xor~14_combout ;
wire \Equal0~15_combout ;
wire \Equal0~16_combout ;
wire \D_ctrl_force_src2_zero~0_combout ;
wire \Equal62~14_combout ;
wire \Equal62~13_combout ;
wire \D_ctrl_force_src2_zero~1_combout ;
wire \Equal62~8_combout ;
wire \D_ctrl_force_src2_zero~2_combout ;
wire \Equal0~13_combout ;
wire \Equal0~2_combout ;
wire \D_ctrl_force_src2_zero~3_combout ;
wire \D_ctrl_force_src2_zero~4_combout ;
wire \Equal62~9_combout ;
wire \D_ctrl_uncond_cti_non_br~1_combout ;
wire \Equal62~10_combout ;
wire \Equal0~3_combout ;
wire \D_op_cmpge~0_combout ;
wire \D_ctrl_exception~13_combout ;
wire \Equal62~11_combout ;
wire \D_op_opx_rsv17~0_combout ;
wire \D_ctrl_exception~14_combout ;
wire \Equal62~2_combout ;
wire \D_op_opx_rsv00~0_combout ;
wire \D_ctrl_exception~15_combout ;
wire \D_ctrl_exception~16_combout ;
wire \D_ctrl_exception~17_combout ;
wire \D_ctrl_exception~18_combout ;
wire \Equal0~12_combout ;
wire \D_ctrl_exception~19_combout ;
wire \Equal62~12_combout ;
wire \Equal62~3_combout ;
wire \Equal62~1_combout ;
wire \D_ctrl_exception~20_combout ;
wire \D_ctrl_exception~23_combout ;
wire \D_ctrl_exception~21_combout ;
wire \Equal0~4_combout ;
wire \D_ctrl_jmp_direct~0_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \D_ctrl_retaddr~2_combout ;
wire \D_ctrl_force_src2_zero~5_combout ;
wire \Equal0~18_combout ;
wire \D_ctrl_force_src2_zero~6_combout ;
wire \D_ctrl_force_src2_zero~7_combout ;
wire \R_ctrl_force_src2_zero~q ;
wire \R_src2_lo[4]~2_combout ;
wire \F_iw[6]~44_combout ;
wire \F_iw[6]~46_combout ;
wire \D_iw[6]~q ;
wire \D_ctrl_src_imm5_shift_rot~0_combout ;
wire \D_ctrl_src_imm5_shift_rot~1_combout ;
wire \R_ctrl_src_imm5_shift_rot~q ;
wire \D_ctrl_implicit_dst_eretaddr~7_combout ;
wire \D_ctrl_unsigned_lo_imm16~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~1_combout ;
wire \Equal0~17_combout ;
wire \D_ctrl_b_is_dst~0_combout ;
wire \D_ctrl_b_is_dst~1_combout ;
wire \D_ctrl_b_is_dst~2_combout ;
wire \R_src2_use_imm~0_combout ;
wire \R_ctrl_br_nxt~0_combout ;
wire \R_ctrl_br_nxt~1_combout ;
wire \R_src2_use_imm~1_combout ;
wire \R_src2_use_imm~q ;
wire \R_src2_lo~3_combout ;
wire \R_src2_lo[0]~8_combout ;
wire \E_src2[0]~q ;
wire \E_shift_rot_cnt[0]~q ;
wire \E_shift_rot_cnt[0]~6 ;
wire \E_shift_rot_cnt[1]~7_combout ;
wire \F_iw[7]~41_combout ;
wire \F_iw[7]~43_combout ;
wire \D_iw[7]~q ;
wire \R_src2_lo[1]~7_combout ;
wire \E_src2[1]~q ;
wire \E_shift_rot_cnt[1]~q ;
wire \E_shift_rot_cnt[1]~8 ;
wire \E_shift_rot_cnt[2]~9_combout ;
wire \R_src2_lo[2]~6_combout ;
wire \E_src2[2]~q ;
wire \E_shift_rot_cnt[2]~q ;
wire \E_stall~0_combout ;
wire \E_shift_rot_cnt[2]~10 ;
wire \E_shift_rot_cnt[3]~11_combout ;
wire \F_iw[9]~35_combout ;
wire \F_iw[9]~37_combout ;
wire \D_iw[9]~q ;
wire \R_src2_lo[3]~5_combout ;
wire \E_src2[3]~q ;
wire \E_shift_rot_cnt[3]~q ;
wire \E_shift_rot_cnt[3]~12 ;
wire \E_shift_rot_cnt[4]~13_combout ;
wire \F_iw[10]~32_combout ;
wire \F_iw[10]~34_combout ;
wire \D_iw[10]~q ;
wire \R_src2_lo[4]~4_combout ;
wire \E_src2[4]~q ;
wire \E_shift_rot_cnt[4]~q ;
wire \E_stall~1_combout ;
wire \E_stall~2_combout ;
wire \D_ctrl_ld_signed~0_combout ;
wire \D_ctrl_ld~2_combout ;
wire \D_ctrl_ld~3_combout ;
wire \R_ctrl_ld~q ;
wire \av_ld_waiting_for_data_nxt~0_combout ;
wire \av_ld_waiting_for_data~q ;
wire \av_ld_waiting_for_data_nxt~1_combout ;
wire \av_ld_aligning_data~q ;
wire \D_ctrl_mem16~0_combout ;
wire \D_ctrl_mem16~1_combout ;
wire \av_ld_align_cycle_nxt[0]~0_combout ;
wire \av_ld_align_cycle[0]~q ;
wire \av_ld_align_cycle_nxt[1]~1_combout ;
wire \av_ld_align_cycle[1]~q ;
wire \av_ld_aligning_data_nxt~0_combout ;
wire \D_ctrl_mem32~0_combout ;
wire \av_ld_aligning_data_nxt~1_combout ;
wire \av_ld_aligning_data_nxt~2_combout ;
wire \E_stall~3_combout ;
wire \E_stall~4_combout ;
wire \E_valid_from_R~3_combout ;
wire \E_valid_from_R~2_combout ;
wire \E_valid_from_R~q ;
wire \D_ctrl_jmp_direct~1_combout ;
wire \R_ctrl_jmp_direct~q ;
wire \R_src1~14_combout ;
wire \E_src1[4]~22_combout ;
wire \F_pc_plus_one[0]~1 ;
wire \F_pc_plus_one[1]~3 ;
wire \F_pc_plus_one[2]~4_combout ;
wire \R_ctrl_br~q ;
wire \D_ctrl_retaddr~3_combout ;
wire \D_ctrl_retaddr~4_combout ;
wire \D_ctrl_retaddr~5_combout ;
wire \Equal0~10_combout ;
wire \D_ctrl_retaddr~6_combout ;
wire \D_ctrl_retaddr~7_combout ;
wire \D_ctrl_retaddr~8_combout ;
wire \R_ctrl_retaddr~q ;
wire \R_src1~15_combout ;
wire \E_src1[4]~q ;
wire \Equal135~0_combout ;
wire \Equal135~1_combout ;
wire \D_op_wrctl~combout ;
wire \R_ctrl_wrctl_inst~q ;
wire \W_ienable_reg_nxt~0_combout ;
wire \W_ienable_reg[4]~q ;
wire \W_ipending_reg_nxt[4]~0_combout ;
wire \W_ipending_reg[4]~q ;
wire \E_src1[3]~23_combout ;
wire \F_pc_plus_one[1]~2_combout ;
wire \E_src1[3]~q ;
wire \W_ienable_reg[3]~q ;
wire \W_ipending_reg_nxt[3]~1_combout ;
wire \W_ipending_reg[3]~q ;
wire \E_src1[2]~24_combout ;
wire \F_pc_plus_one[0]~0_combout ;
wire \E_src1[2]~q ;
wire \W_ienable_reg[2]~q ;
wire \W_ipending_reg_nxt[2]~2_combout ;
wire \W_ipending_reg[2]~q ;
wire \R_src1[1]~16_combout ;
wire \E_src1[1]~q ;
wire \W_ienable_reg[1]~q ;
wire \W_ipending_reg_nxt[1]~3_combout ;
wire \W_ipending_reg[1]~q ;
wire \D_iw[1]~0_combout ;
wire \R_src1[0]~17_combout ;
wire \E_src1[0]~q ;
wire \W_ienable_reg[0]~q ;
wire \W_ipending_reg_nxt[0]~4_combout ;
wire \W_ipending_reg[0]~q ;
wire \E_wrctl_estatus~0_combout ;
wire \E_wrctl_status~1_combout ;
wire \W_estatus_reg_inst_nxt~0_combout ;
wire \D_ctrl_exception~7_combout ;
wire \D_ctrl_exception~24_combout ;
wire \D_ctrl_exception~10_combout ;
wire \D_ctrl_exception~11_combout ;
wire \D_ctrl_exception~12_combout ;
wire \D_ctrl_implicit_dst_eretaddr~0_combout ;
wire \D_ctrl_implicit_dst_eretaddr~1_combout ;
wire \D_ctrl_implicit_dst_eretaddr~2_combout ;
wire \D_ctrl_exception~22_combout ;
wire \R_ctrl_exception~q ;
wire \W_estatus_reg_inst_nxt~1_combout ;
wire \W_estatus_reg~q ;
wire \E_wrctl_bstatus~0_combout ;
wire \D_ctrl_break~0_combout ;
wire \R_ctrl_break~q ;
wire \W_bstatus_reg_inst_nxt~0_combout ;
wire \W_bstatus_reg_inst_nxt~1_combout ;
wire \W_bstatus_reg~q ;
wire \E_wrctl_status~0_combout ;
wire \W_status_reg_pie_inst_nxt~0_combout ;
wire \W_status_reg_pie_inst_nxt~1_combout ;
wire \D_op_eret~combout ;
wire \F_pc_sel_nxt.10~0_combout ;
wire \W_status_reg_pie_inst_nxt~2_combout ;
wire \W_status_reg_pie~q ;
wire \D_iw[1]~1_combout ;
wire \D_iw[1]~2_combout ;
wire \F_iw[11]~17_combout ;
wire \D_iw[11]~q ;
wire \Equal62~0_combout ;
wire \Equal0~5_combout ;
wire \D_ctrl_alu_subtract~8_combout ;
wire \D_ctrl_alu_subtract~9_combout ;
wire \D_ctrl_alu_subtract~5_combout ;
wire \D_ctrl_alu_subtract~10_combout ;
wire \E_alu_sub~0_combout ;
wire \E_alu_sub~q ;
wire \E_src2[5]~15_combout ;
wire \R_src2_lo[6]~0_combout ;
wire \E_src2[6]~q ;
wire \Add1~0_combout ;
wire \E_src1[6]~20_combout ;
wire \F_pc_plus_one[2]~5 ;
wire \F_pc_plus_one[3]~7 ;
wire \F_pc_plus_one[4]~8_combout ;
wire \E_src1[6]~q ;
wire \R_src2_lo[5]~1_combout ;
wire \E_src2[5]~q ;
wire \Add1~1_combout ;
wire \E_src1[5]~21_combout ;
wire \F_pc_plus_one[3]~6_combout ;
wire \E_src1[5]~q ;
wire \Add1~2_combout ;
wire \Add1~3_combout ;
wire \Add1~4_combout ;
wire \Add1~5_combout ;
wire \Add1~6_combout ;
wire \Add1~8_cout ;
wire \Add1~10 ;
wire \Add1~12 ;
wire \Add1~14 ;
wire \Add1~16 ;
wire \Add1~18 ;
wire \Add1~20 ;
wire \Add1~21_combout ;
wire \D_logic_op_raw[1]~0_combout ;
wire \D_ctrl_alu_force_xor~10_combout ;
wire \D_ctrl_alu_force_xor~11_combout ;
wire \D_ctrl_alu_force_xor~13_combout ;
wire \D_ctrl_alu_force_xor~12_combout ;
wire \D_logic_op[1]~0_combout ;
wire \R_logic_op[1]~q ;
wire \D_logic_op[0]~1_combout ;
wire \R_logic_op[0]~q ;
wire \E_logic_result[6]~0_combout ;
wire \Equal0~9_combout ;
wire \Equal0~11_combout ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_logic~combout ;
wire \R_ctrl_logic~q ;
wire \W_alu_result[6]~20_combout ;
wire \D_ctrl_shift_rot_right~0_combout ;
wire \D_ctrl_shift_rot_right~1_combout ;
wire \R_ctrl_shift_rot_right~q ;
wire \E_shift_rot_result_nxt[5]~18_combout ;
wire \E_shift_rot_result[5]~q ;
wire \E_shift_rot_result_nxt[4]~22_combout ;
wire \E_shift_rot_result[4]~q ;
wire \E_shift_rot_result_nxt[3]~23_combout ;
wire \E_shift_rot_result[3]~q ;
wire \E_shift_rot_result_nxt[2]~24_combout ;
wire \E_shift_rot_result[2]~q ;
wire \E_shift_rot_result_nxt[1]~26_combout ;
wire \E_shift_rot_result[1]~q ;
wire \E_shift_rot_result_nxt[0]~28_combout ;
wire \E_shift_rot_result[0]~q ;
wire \R_ctrl_rot_right_nxt~0_combout ;
wire \R_ctrl_rot_right~q ;
wire \D_ctrl_shift_logical~1_combout ;
wire \D_ctrl_shift_logical~2_combout ;
wire \R_ctrl_shift_logical~q ;
wire \E_shift_rot_fill_bit~0_combout ;
wire \E_shift_rot_result_nxt[31]~30_combout ;
wire \R_src1[31]~18_combout ;
wire \E_src1[31]~q ;
wire \E_shift_rot_result[31]~q ;
wire \E_shift_rot_result_nxt[30]~31_combout ;
wire \R_src1[30]~19_combout ;
wire \E_src1[30]~q ;
wire \E_shift_rot_result[30]~q ;
wire \E_shift_rot_result_nxt[29]~29_combout ;
wire \R_src1[29]~20_combout ;
wire \E_src1[29]~q ;
wire \E_shift_rot_result[29]~q ;
wire \E_shift_rot_result_nxt[28]~27_combout ;
wire \R_src1[28]~21_combout ;
wire \E_src1[28]~q ;
wire \E_shift_rot_result[28]~q ;
wire \E_shift_rot_result_nxt[27]~25_combout ;
wire \R_src1[27]~22_combout ;
wire \E_src1[27]~q ;
wire \E_shift_rot_result[27]~q ;
wire \E_shift_rot_result_nxt[26]~1_combout ;
wire \F_iw[30]~49_combout ;
wire \F_iw[30]~50_combout ;
wire \D_iw[30]~q ;
wire \E_src1[26]~0_combout ;
wire \F_pc_plus_one[4]~9 ;
wire \F_pc_plus_one[5]~11 ;
wire \F_pc_plus_one[6]~13 ;
wire \F_pc_plus_one[7]~15 ;
wire \F_pc_plus_one[8]~17 ;
wire \F_pc_plus_one[9]~19 ;
wire \F_pc_plus_one[10]~21 ;
wire \F_pc_plus_one[11]~23 ;
wire \F_pc_plus_one[12]~25 ;
wire \F_pc_plus_one[13]~27 ;
wire \F_pc_plus_one[14]~29 ;
wire \F_pc_plus_one[15]~31 ;
wire \F_pc_plus_one[16]~33 ;
wire \F_pc_plus_one[17]~35 ;
wire \F_pc_plus_one[18]~37 ;
wire \F_pc_plus_one[19]~39 ;
wire \F_pc_plus_one[20]~41 ;
wire \F_pc_plus_one[21]~43 ;
wire \F_pc_plus_one[22]~45 ;
wire \F_pc_plus_one[23]~47 ;
wire \F_pc_plus_one[24]~48_combout ;
wire \E_src1[26]~q ;
wire \E_shift_rot_result[26]~q ;
wire \E_shift_rot_result_nxt[25]~2_combout ;
wire \F_iw[29]~51_combout ;
wire \F_iw[29]~52_combout ;
wire \D_iw[29]~q ;
wire \E_src1[25]~1_combout ;
wire \F_pc_plus_one[23]~46_combout ;
wire \E_src1[25]~q ;
wire \E_shift_rot_result[25]~q ;
wire \E_shift_rot_result_nxt[24]~3_combout ;
wire \F_iw[28]~53_combout ;
wire \F_iw[28]~54_combout ;
wire \D_iw[28]~q ;
wire \E_src1[24]~2_combout ;
wire \F_pc_plus_one[22]~44_combout ;
wire \E_src1[24]~q ;
wire \E_shift_rot_result[24]~q ;
wire \E_shift_rot_result_nxt[23]~4_combout ;
wire \F_iw[27]~55_combout ;
wire \F_iw[27]~56_combout ;
wire \D_iw[27]~q ;
wire \E_src1[23]~3_combout ;
wire \F_pc_plus_one[21]~42_combout ;
wire \E_src1[23]~q ;
wire \E_shift_rot_result[23]~q ;
wire \E_shift_rot_result_nxt[22]~5_combout ;
wire \F_iw[26]~57_combout ;
wire \F_iw[26]~58_combout ;
wire \D_iw[26]~q ;
wire \E_src1[22]~4_combout ;
wire \F_pc_plus_one[20]~40_combout ;
wire \E_src1[22]~q ;
wire \E_shift_rot_result[22]~q ;
wire \E_shift_rot_result_nxt[21]~6_combout ;
wire \F_iw[25]~59_combout ;
wire \F_iw[25]~60_combout ;
wire \D_iw[25]~q ;
wire \E_src1[21]~5_combout ;
wire \F_pc_plus_one[19]~38_combout ;
wire \E_src1[21]~q ;
wire \E_shift_rot_result[21]~q ;
wire \E_shift_rot_result_nxt[20]~7_combout ;
wire \F_iw[24]~61_combout ;
wire \F_iw[24]~62_combout ;
wire \D_iw[24]~q ;
wire \E_src1[20]~6_combout ;
wire \F_pc_plus_one[18]~36_combout ;
wire \E_src1[20]~q ;
wire \E_shift_rot_result[20]~q ;
wire \E_shift_rot_result_nxt[19]~8_combout ;
wire \F_iw[23]~63_combout ;
wire \F_iw[23]~64_combout ;
wire \D_iw[23]~q ;
wire \E_src1[19]~7_combout ;
wire \F_pc_plus_one[17]~34_combout ;
wire \E_src1[19]~q ;
wire \E_shift_rot_result[19]~q ;
wire \E_shift_rot_result_nxt[18]~9_combout ;
wire \F_iw[22]~65_combout ;
wire \F_iw[22]~66_combout ;
wire \D_iw[22]~q ;
wire \E_src1[18]~8_combout ;
wire \F_pc_plus_one[16]~32_combout ;
wire \E_src1[18]~q ;
wire \E_shift_rot_result[18]~q ;
wire \E_shift_rot_result_nxt[17]~10_combout ;
wire \F_iw[21]~47_combout ;
wire \F_iw[21]~48_combout ;
wire \D_iw[21]~q ;
wire \E_src1[17]~9_combout ;
wire \F_pc_plus_one[15]~30_combout ;
wire \E_src1[17]~q ;
wire \E_shift_rot_result[17]~q ;
wire \E_shift_rot_result_nxt[16]~11_combout ;
wire \F_iw[20]~67_combout ;
wire \F_iw[20]~68_combout ;
wire \D_iw[20]~q ;
wire \E_src1[16]~10_combout ;
wire \F_pc_plus_one[14]~28_combout ;
wire \E_src1[16]~q ;
wire \E_shift_rot_result[16]~q ;
wire \E_shift_rot_result_nxt[15]~12_combout ;
wire \F_iw[19]~69_combout ;
wire \F_iw[19]~70_combout ;
wire \D_iw[19]~q ;
wire \E_src1[15]~11_combout ;
wire \F_pc_plus_one[13]~26_combout ;
wire \E_src1[15]~q ;
wire \E_shift_rot_result[15]~q ;
wire \E_shift_rot_result_nxt[14]~13_combout ;
wire \F_iw[18]~71_combout ;
wire \F_iw[18]~72_combout ;
wire \F_iw[18]~73_combout ;
wire \D_iw[18]~q ;
wire \E_src1[14]~12_combout ;
wire \F_pc_plus_one[12]~24_combout ;
wire \E_src1[14]~q ;
wire \E_shift_rot_result[14]~q ;
wire \E_shift_rot_result_nxt[13]~14_combout ;
wire \F_iw[17]~74_combout ;
wire \F_iw[17]~75_combout ;
wire \F_iw[17]~79_combout ;
wire \D_iw[17]~q ;
wire \E_src1[13]~13_combout ;
wire \F_pc_plus_one[11]~22_combout ;
wire \E_src1[13]~q ;
wire \E_shift_rot_result[13]~q ;
wire \E_shift_rot_result_nxt[12]~15_combout ;
wire \E_src1[12]~14_combout ;
wire \F_pc_plus_one[10]~20_combout ;
wire \E_src1[12]~q ;
wire \E_shift_rot_result[12]~q ;
wire \E_shift_rot_result_nxt[11]~16_combout ;
wire \E_src1[11]~15_combout ;
wire \F_pc_plus_one[9]~18_combout ;
wire \E_src1[11]~q ;
wire \E_shift_rot_result[11]~q ;
wire \E_shift_rot_result_nxt[10]~17_combout ;
wire \E_src1[10]~16_combout ;
wire \F_pc_plus_one[8]~16_combout ;
wire \E_src1[10]~q ;
wire \E_shift_rot_result[10]~q ;
wire \E_shift_rot_result_nxt[9]~20_combout ;
wire \E_src1[9]~17_combout ;
wire \F_pc_plus_one[7]~14_combout ;
wire \E_src1[9]~q ;
wire \E_shift_rot_result[9]~q ;
wire \E_shift_rot_result_nxt[8]~21_combout ;
wire \E_src1[8]~18_combout ;
wire \F_pc_plus_one[6]~12_combout ;
wire \E_src1[8]~q ;
wire \E_shift_rot_result[8]~q ;
wire \E_shift_rot_result_nxt[7]~19_combout ;
wire \E_src1[7]~19_combout ;
wire \F_pc_plus_one[5]~10_combout ;
wire \E_src1[7]~q ;
wire \E_shift_rot_result[7]~q ;
wire \E_shift_rot_result_nxt[6]~0_combout ;
wire \E_shift_rot_result[6]~q ;
wire \D_op_rdctl~combout ;
wire \R_ctrl_rd_ctl_reg~q ;
wire \Equal0~6_combout ;
wire \D_ctrl_br_cmp~2_combout ;
wire \D_ctrl_br_cmp~5_combout ;
wire \D_ctrl_br_cmp~3_combout ;
wire \D_ctrl_br_cmp~4_combout ;
wire \R_ctrl_br_cmp~q ;
wire \E_alu_result~0_combout ;
wire \E_src2[26]~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~2_combout ;
wire \D_ctrl_unsigned_lo_imm16~3_combout ;
wire \R_ctrl_unsigned_lo_imm16~q ;
wire \R_src2_hi~0_combout ;
wire \E_src2[26]~q ;
wire \Add1~23_combout ;
wire \E_src2[25]~1_combout ;
wire \E_src2[25]~q ;
wire \Add1~24_combout ;
wire \E_src2[24]~2_combout ;
wire \E_src2[24]~q ;
wire \Add1~25_combout ;
wire \E_src2[23]~3_combout ;
wire \E_src2[23]~q ;
wire \Add1~26_combout ;
wire \E_src2[22]~4_combout ;
wire \E_src2[22]~q ;
wire \Add1~27_combout ;
wire \E_src2[21]~5_combout ;
wire \E_src2[21]~q ;
wire \Add1~28_combout ;
wire \E_src2[20]~6_combout ;
wire \E_src2[20]~q ;
wire \Add1~29_combout ;
wire \E_src2[19]~7_combout ;
wire \E_src2[19]~q ;
wire \Add1~30_combout ;
wire \E_src2[18]~8_combout ;
wire \E_src2[18]~q ;
wire \Add1~31_combout ;
wire \E_src2[17]~9_combout ;
wire \E_src2[17]~q ;
wire \Add1~32_combout ;
wire \E_src2[16]~10_combout ;
wire \E_src2[16]~q ;
wire \Add1~33_combout ;
wire \R_src2_lo[15]~9_combout ;
wire \E_src2[15]~q ;
wire \Add1~34_combout ;
wire \R_src2_lo[14]~10_combout ;
wire \E_src2[14]~q ;
wire \Add1~35_combout ;
wire \R_src2_lo[13]~11_combout ;
wire \E_src2[13]~q ;
wire \Add1~36_combout ;
wire \R_src2_lo[12]~12_combout ;
wire \E_src2[12]~q ;
wire \Add1~37_combout ;
wire \R_src2_lo[11]~13_combout ;
wire \E_src2[11]~q ;
wire \Add1~38_combout ;
wire \R_src2_lo[10]~14_combout ;
wire \E_src2[10]~q ;
wire \Add1~39_combout ;
wire \R_src2_lo[9]~15_combout ;
wire \E_src2[9]~q ;
wire \Add1~40_combout ;
wire \R_src2_lo[8]~16_combout ;
wire \E_src2[8]~q ;
wire \Add1~41_combout ;
wire \R_src2_lo[7]~17_combout ;
wire \E_src2[7]~q ;
wire \Add1~42_combout ;
wire \Add1~22 ;
wire \Add1~44 ;
wire \Add1~46 ;
wire \Add1~48 ;
wire \Add1~50 ;
wire \Add1~52 ;
wire \Add1~54 ;
wire \Add1~56 ;
wire \Add1~58 ;
wire \Add1~60 ;
wire \Add1~62 ;
wire \Add1~64 ;
wire \Add1~66 ;
wire \Add1~68 ;
wire \Add1~70 ;
wire \Add1~72 ;
wire \Add1~74 ;
wire \Add1~76 ;
wire \Add1~78 ;
wire \Add1~80 ;
wire \Add1~81_combout ;
wire \E_logic_result[26]~1_combout ;
wire \W_alu_result[26]~0_combout ;
wire \Add1~79_combout ;
wire \E_logic_result[25]~2_combout ;
wire \W_alu_result[25]~1_combout ;
wire \Add1~77_combout ;
wire \E_logic_result[24]~3_combout ;
wire \W_alu_result[24]~2_combout ;
wire \Add1~75_combout ;
wire \E_logic_result[23]~4_combout ;
wire \W_alu_result[23]~3_combout ;
wire \Add1~73_combout ;
wire \E_logic_result[22]~5_combout ;
wire \W_alu_result[22]~4_combout ;
wire \Add1~71_combout ;
wire \E_logic_result[21]~6_combout ;
wire \W_alu_result[21]~5_combout ;
wire \Add1~69_combout ;
wire \E_logic_result[20]~7_combout ;
wire \W_alu_result[20]~6_combout ;
wire \Add1~67_combout ;
wire \E_logic_result[19]~8_combout ;
wire \W_alu_result[19]~7_combout ;
wire \Add1~65_combout ;
wire \E_logic_result[18]~9_combout ;
wire \W_alu_result[18]~8_combout ;
wire \Add1~63_combout ;
wire \E_logic_result[17]~10_combout ;
wire \W_alu_result[17]~9_combout ;
wire \Add1~61_combout ;
wire \E_logic_result[16]~11_combout ;
wire \W_alu_result[16]~10_combout ;
wire \Add1~59_combout ;
wire \E_logic_result[15]~12_combout ;
wire \W_alu_result[15]~11_combout ;
wire \Add1~57_combout ;
wire \E_logic_result[14]~13_combout ;
wire \W_alu_result[14]~12_combout ;
wire \Add1~55_combout ;
wire \E_logic_result[13]~14_combout ;
wire \W_alu_result[13]~13_combout ;
wire \Add1~53_combout ;
wire \E_logic_result[12]~15_combout ;
wire \W_alu_result[12]~14_combout ;
wire \Add1~51_combout ;
wire \E_logic_result[11]~16_combout ;
wire \W_alu_result[11]~15_combout ;
wire \Add1~49_combout ;
wire \E_logic_result[10]~17_combout ;
wire \W_alu_result[10]~16_combout ;
wire \Add1~19_combout ;
wire \E_logic_result[5]~18_combout ;
wire \W_alu_result[5]~21_combout ;
wire \Add1~43_combout ;
wire \E_logic_result[7]~19_combout ;
wire \W_alu_result[7]~19_combout ;
wire \Add1~47_combout ;
wire \E_logic_result[9]~20_combout ;
wire \W_alu_result[9]~17_combout ;
wire \Add1~45_combout ;
wire \E_logic_result[8]~21_combout ;
wire \W_alu_result[8]~18_combout ;
wire \Add1~17_combout ;
wire \E_logic_result[4]~22_combout ;
wire \W_alu_result[4]~22_combout ;
wire \Add1~15_combout ;
wire \E_logic_result[3]~23_combout ;
wire \W_alu_result[3]~23_combout ;
wire \Add1~13_combout ;
wire \E_logic_result[2]~24_combout ;
wire \W_alu_result[2]~24_combout ;
wire \d_writedata[24]~0_combout ;
wire \D_ctrl_mem8~0_combout ;
wire \D_ctrl_mem8~1_combout ;
wire \d_writedata[25]~1_combout ;
wire \d_writedata[26]~2_combout ;
wire \d_writedata[27]~3_combout ;
wire \d_writedata[28]~4_combout ;
wire \d_writedata[29]~5_combout ;
wire \d_writedata[30]~6_combout ;
wire \d_writedata[31]~7_combout ;
wire \d_read_nxt~combout ;
wire \E_st_stall~combout ;
wire \Add1~9_combout ;
wire \Add1~11_combout ;
wire \E_mem_byte_en[0]~0_combout ;
wire \E_mem_byte_en[1]~1_combout ;
wire \i_read_nxt~0_combout ;
wire \D_ctrl_uncond_cti_non_br~0_combout ;
wire \D_ctrl_uncond_cti_non_br~2_combout ;
wire \R_ctrl_uncond_cti_non_br~q ;
wire \Equal0~20_combout ;
wire \R_ctrl_br_uncond~q ;
wire \R_compare_op[1]~q ;
wire \D_logic_op_raw[0]~1_combout ;
wire \R_compare_op[0]~q ;
wire \Equal127~0_combout ;
wire \Equal127~1_combout ;
wire \Equal127~2_combout ;
wire \Equal127~3_combout ;
wire \Equal127~4_combout ;
wire \Equal127~5_combout ;
wire \Equal127~6_combout ;
wire \R_src2_hi[15]~1_combout ;
wire \R_src2_hi[15]~2_combout ;
wire \E_src2[31]~q ;
wire \E_logic_result[31]~25_combout ;
wire \E_src2[30]~11_combout ;
wire \E_src2[30]~q ;
wire \E_logic_result[30]~26_combout ;
wire \E_src2[29]~12_combout ;
wire \E_src2[29]~q ;
wire \E_logic_result[29]~27_combout ;
wire \Equal127~7_combout ;
wire \E_src2[28]~13_combout ;
wire \E_src2[28]~q ;
wire \E_logic_result[28]~28_combout ;
wire \E_src2[27]~14_combout ;
wire \E_src2[27]~q ;
wire \E_logic_result[27]~29_combout ;
wire \E_logic_result[1]~30_combout ;
wire \E_logic_result[0]~31_combout ;
wire \Equal127~8_combout ;
wire \Equal127~9_combout ;
wire \E_cmp_result~0_combout ;
wire \E_invert_arith_src_msb~0_combout ;
wire \E_invert_arith_src_msb~1_combout ;
wire \E_invert_arith_src_msb~q ;
wire \Add1~83_combout ;
wire \E_arith_src1[31]~combout ;
wire \Add1~84_combout ;
wire \Add1~85_combout ;
wire \Add1~86_combout ;
wire \Add1~87_combout ;
wire \Add1~82 ;
wire \Add1~89 ;
wire \Add1~91 ;
wire \Add1~93 ;
wire \Add1~95 ;
wire \Add1~97 ;
wire \Add1~98_combout ;
wire \E_cmp_result~1_combout ;
wire \W_cmp_result~q ;
wire \F_pc_sel_nxt~0_combout ;
wire \F_pc_no_crst_nxt[24]~0_combout ;
wire \F_pc_no_crst_nxt[24]~1_combout ;
wire \F_pc_no_crst_nxt[23]~2_combout ;
wire \F_pc_no_crst_nxt[23]~3_combout ;
wire \F_pc_no_crst_nxt[22]~4_combout ;
wire \F_pc_no_crst_nxt[21]~5_combout ;
wire \F_pc_no_crst_nxt[20]~6_combout ;
wire \F_pc_no_crst_nxt[19]~7_combout ;
wire \F_pc_no_crst_nxt[18]~8_combout ;
wire \F_pc_no_crst_nxt[17]~9_combout ;
wire \F_pc_no_crst_nxt[16]~10_combout ;
wire \F_pc_no_crst_nxt[15]~11_combout ;
wire \F_pc_no_crst_nxt[14]~12_combout ;
wire \F_pc_no_crst_nxt[13]~13_combout ;
wire \F_pc_no_crst_nxt[12]~14_combout ;
wire \F_pc_no_crst_nxt[11]~15_combout ;
wire \F_pc_no_crst_nxt[10]~16_combout ;
wire \F_pc_no_crst_nxt[10]~17_combout ;
wire \F_pc_no_crst_nxt[8]~18_combout ;
wire \F_pc_no_crst_nxt[9]~19_combout ;
wire \F_pc_no_crst_nxt[9]~20_combout ;
wire \F_pc_no_crst_nxt[0]~21_combout ;
wire \F_pc_no_crst_nxt[1]~22_combout ;
wire \F_pc_no_crst_nxt[2]~23_combout ;
wire \F_pc_no_crst_nxt[3]~24_combout ;
wire \F_pc_no_crst_nxt[4]~25_combout ;
wire \F_pc_no_crst_nxt[5]~26_combout ;
wire \F_pc_no_crst_nxt[6]~27_combout ;
wire \F_pc_no_crst_nxt[7]~28_combout ;
wire \E_st_data[10]~0_combout ;
wire \E_mem_byte_en[2]~2_combout ;
wire \E_mem_byte_en[3]~3_combout ;
wire \hbreak_enabled~0_combout ;
wire \E_st_data[8]~1_combout ;
wire \E_st_data[9]~2_combout ;
wire \E_st_data[11]~3_combout ;
wire \E_st_data[12]~4_combout ;
wire \E_st_data[13]~5_combout ;
wire \E_st_data[14]~6_combout ;
wire \E_st_data[15]~7_combout ;
wire \d_byteenable[3]~0_combout ;
wire \E_st_data[16]~8_combout ;
wire \E_st_data[17]~9_combout ;
wire \E_st_data[18]~10_combout ;
wire \E_st_data[19]~11_combout ;
wire \E_st_data[20]~12_combout ;
wire \E_st_data[21]~13_combout ;
wire \E_st_data[22]~14_combout ;
wire \E_st_data[23]~15_combout ;


niosII_niosII_cpu_cpu_nios2_oci the_niosII_cpu_cpu_nios2_oci(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.sr_0(sr_0),
	.jtag_break(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_oci_debug|jtag_break~q ),
	.readdata_4(readdata_4),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.r_sync_rst(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.hbreak_enabled(hbreak_enabled1),
	.WideOr1(WideOr11),
	.rf_source_valid(rf_source_valid),
	.uav_write(uav_write),
	.r_early_rst(r_early_rst),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_411,src_data_40,src_data_39,src_data_38}),
	.oci_ienable_4(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[4]~q ),
	.oci_ienable_3(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[3]~q ),
	.oci_ienable_2(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[2]~q ),
	.oci_ienable_1(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.oci_ienable_0(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.oci_single_step_mode(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.readdata_0(readdata_0),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.readdata_3(readdata_3),
	.debugaccess_nxt(src_payload1),
	.writedata_nxt({src_payload42,src_payload29,src_payload30,src_payload31,src_payload32,src_payload33,src_payload34,src_payload35,src_payload36,src_payload37,src_payload28,src_payload38,src_payload39,src_payload40,src_payload41,src_payload18,src_payload22,src_payload21,src_payload17,
src_payload19,src_payload16,src_payload23,src_payload24,src_payload25,src_payload26,src_payload27,src_payload20,src_payload13,src_payload14,src_payload15,src_payload12,src_payload2}),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.readdata_11(readdata_11),
	.readdata_13(readdata_13),
	.readdata_16(readdata_16),
	.readdata_12(readdata_12),
	.readdata_5(readdata_5),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_10(readdata_10),
	.readdata_9(readdata_9),
	.readdata_8(readdata_8),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.readdata_21(readdata_21),
	.readdata_30(readdata_30),
	.readdata_29(readdata_29),
	.readdata_28(readdata_28),
	.readdata_27(readdata_27),
	.readdata_26(readdata_261),
	.readdata_25(readdata_251),
	.readdata_24(readdata_241),
	.readdata_23(readdata_23),
	.readdata_22(readdata_22),
	.readdata_20(readdata_20),
	.readdata_19(readdata_19),
	.readdata_18(readdata_18),
	.readdata_17(readdata_17),
	.readdata_31(readdata_311),
	.resetrequest(debug_reset_request),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

niosII_niosII_cpu_cpu_register_bank_b_module niosII_cpu_cpu_register_bank_b(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.q_b_0(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_7(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_26(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_24(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_16(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_27(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_28(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_29(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_30(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_31(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.D_iw_26(\D_iw[26]~q ),
	.D_iw_25(\D_iw[25]~q ),
	.D_iw_24(\D_iw[24]~q ),
	.D_iw_23(\D_iw[23]~q ),
	.D_iw_22(\D_iw[22]~q ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~4_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~6_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~8_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~10_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~11_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~12_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~13_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~14_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~15_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~16_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~17_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~18_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~19_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~20_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~21_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~22_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~23_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~24_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~25_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~26_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~27_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~28_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~29_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~30_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~31_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~32_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~33_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~34_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~35_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~36_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~37_combout ));

niosII_niosII_cpu_cpu_register_bank_a_module niosII_cpu_cpu_register_bank_a(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.q_b_6(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_5(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_3(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_2(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_1(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_26(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_24(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_16(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_31(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_30(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_29(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_28(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.D_iw_30(\D_iw[30]~q ),
	.D_iw_29(\D_iw[29]~q ),
	.D_iw_28(\D_iw[28]~q ),
	.D_iw_27(\D_iw[27]~q ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~4_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~6_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~8_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~10_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~11_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~12_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~13_combout ),
	.D_iw_31(\D_iw[31]~q ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~14_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~15_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~16_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~17_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~18_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~19_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~20_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~21_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~22_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~23_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~24_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~25_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~26_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~27_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~28_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~29_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~30_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~31_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~32_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~33_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~34_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~35_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~36_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~37_combout ));

dffeas \W_alu_result[0] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[0]~25_combout ),
	.asdata(\E_shift_rot_result[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[0]~q ),
	.prn(vcc));
defparam \W_alu_result[0] .is_wysiwyg = "true";
defparam \W_alu_result[0] .power_up = "low";

dffeas \W_alu_result[1] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[1]~26_combout ),
	.asdata(\E_shift_rot_result[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[1]~q ),
	.prn(vcc));
defparam \W_alu_result[1] .is_wysiwyg = "true";
defparam \W_alu_result[1] .power_up = "low";

cycloneive_lcell_comb \Add1~88 (
	.dataa(\Add1~87_combout ),
	.datab(\E_src1[27]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~82 ),
	.combout(\Add1~88_combout ),
	.cout(\Add1~89 ));
defparam \Add1~88 .lut_mask = 16'h96EF;
defparam \Add1~88 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~90 (
	.dataa(\Add1~86_combout ),
	.datab(\E_src1[28]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~89 ),
	.combout(\Add1~90_combout ),
	.cout(\Add1~91 ));
defparam \Add1~90 .lut_mask = 16'h967F;
defparam \Add1~90 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~92 (
	.dataa(\Add1~85_combout ),
	.datab(\E_src1[29]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~91 ),
	.combout(\Add1~92_combout ),
	.cout(\Add1~93 ));
defparam \Add1~92 .lut_mask = 16'h96EF;
defparam \Add1~92 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~94 (
	.dataa(\Add1~84_combout ),
	.datab(\E_src1[30]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~93 ),
	.combout(\Add1~94_combout ),
	.cout(\Add1~95 ));
defparam \Add1~94 .lut_mask = 16'h967F;
defparam \Add1~94 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~96 (
	.dataa(\Add1~83_combout ),
	.datab(\E_arith_src1[31]~combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~95 ),
	.combout(\Add1~96_combout ),
	.cout(\Add1~97 ));
defparam \Add1~96 .lut_mask = 16'h96EF;
defparam \Add1~96 .sum_lutc_input = "cin";

dffeas \av_ld_byte2_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte2_data[7]~0_combout ),
	.asdata(\av_ld_byte3_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[7] .power_up = "low";

dffeas \av_ld_byte2_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte2_data[6]~1_combout ),
	.asdata(\av_ld_byte3_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[6] .power_up = "low";

dffeas \av_ld_byte2_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte2_data[5]~2_combout ),
	.asdata(\av_ld_byte3_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[5] .power_up = "low";

dffeas \av_ld_byte2_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte2_data[4]~3_combout ),
	.asdata(\av_ld_byte3_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[4] .power_up = "low";

dffeas \av_ld_byte2_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte2_data[3]~4_combout ),
	.asdata(\av_ld_byte3_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[3] .power_up = "low";

dffeas \av_ld_byte2_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte2_data[2]~5_combout ),
	.asdata(\av_ld_byte3_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[2] .power_up = "low";

dffeas \av_ld_byte2_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte2_data[1]~6_combout ),
	.asdata(\av_ld_byte3_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[1] .power_up = "low";

dffeas \av_ld_byte2_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte2_data[0]~7_combout ),
	.asdata(\av_ld_byte3_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[0] .power_up = "low";

dffeas \av_ld_byte1_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte1_data[7]~0_combout ),
	.asdata(\av_ld_byte2_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[7] .power_up = "low";

dffeas \av_ld_byte1_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte1_data[6]~1_combout ),
	.asdata(\av_ld_byte2_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[6] .power_up = "low";

dffeas \av_ld_byte1_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte1_data[5]~2_combout ),
	.asdata(\av_ld_byte2_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[5] .power_up = "low";

dffeas \av_ld_byte1_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte1_data[4]~3_combout ),
	.asdata(\av_ld_byte2_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[4] .power_up = "low";

dffeas \av_ld_byte1_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte1_data[3]~4_combout ),
	.asdata(\av_ld_byte2_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[3] .power_up = "low";

dffeas \av_ld_byte1_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte1_data[2]~5_combout ),
	.asdata(\av_ld_byte2_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[2] .power_up = "low";

dffeas \av_ld_byte1_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte1_data[1]~6_combout ),
	.asdata(\av_ld_byte2_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[1] .power_up = "low";

dffeas \av_ld_byte1_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte1_data[0]~7_combout ),
	.asdata(\av_ld_byte2_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[0] .power_up = "low";

cycloneive_lcell_comb \W_alu_result[0]~25 (
	.dataa(\Add1~9_combout ),
	.datab(\E_logic_result[0]~31_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[0]~25_combout ),
	.cout());
defparam \W_alu_result[0]~25 .lut_mask = 16'hAACC;
defparam \W_alu_result[0]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[1]~26 (
	.dataa(\Add1~11_combout ),
	.datab(\E_logic_result[1]~30_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[1]~26_combout ),
	.cout());
defparam \W_alu_result[1]~26 .lut_mask = 16'hAACC;
defparam \W_alu_result[1]~26 .sum_lutc_input = "datac";

dffeas \W_alu_result[27] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[27]~27_combout ),
	.asdata(\E_shift_rot_result[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[27]~q ),
	.prn(vcc));
defparam \W_alu_result[27] .is_wysiwyg = "true";
defparam \W_alu_result[27] .power_up = "low";

dffeas \W_alu_result[28] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[28]~28_combout ),
	.asdata(\E_shift_rot_result[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[28]~q ),
	.prn(vcc));
defparam \W_alu_result[28] .is_wysiwyg = "true";
defparam \W_alu_result[28] .power_up = "low";

dffeas \W_alu_result[29] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[29]~29_combout ),
	.asdata(\E_shift_rot_result[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[29]~q ),
	.prn(vcc));
defparam \W_alu_result[29] .is_wysiwyg = "true";
defparam \W_alu_result[29] .power_up = "low";

dffeas \W_alu_result[30] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[30]~30_combout ),
	.asdata(\E_shift_rot_result[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[30]~q ),
	.prn(vcc));
defparam \W_alu_result[30] .is_wysiwyg = "true";
defparam \W_alu_result[30] .power_up = "low";

dffeas \W_alu_result[31] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[31]~31_combout ),
	.asdata(\E_shift_rot_result[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[31]~q ),
	.prn(vcc));
defparam \W_alu_result[31] .is_wysiwyg = "true";
defparam \W_alu_result[31] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte2_data[7]~0 (
	.dataa(src_payload4),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[7]~0_combout ),
	.cout());
defparam \av_ld_byte2_data[7]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[7]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[6]~1 (
	.dataa(src_payload5),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[6]~1_combout ),
	.cout());
defparam \av_ld_byte2_data[6]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[6]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[5]~2 (
	.dataa(src_payload6),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[5]~2_combout ),
	.cout());
defparam \av_ld_byte2_data[5]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[5]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[4]~3 (
	.dataa(src_payload7),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[4]~3_combout ),
	.cout());
defparam \av_ld_byte2_data[4]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[4]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[3]~4 (
	.dataa(src_payload8),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[3]~4_combout ),
	.cout());
defparam \av_ld_byte2_data[3]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[2]~5 (
	.dataa(src_payload9),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[2]~5_combout ),
	.cout());
defparam \av_ld_byte2_data[2]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[1]~6 (
	.dataa(src_payload10),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[1]~6_combout ),
	.cout());
defparam \av_ld_byte2_data[1]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[1]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[0]~7 (
	.dataa(src_payload11),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[0]~7_combout ),
	.cout());
defparam \av_ld_byte2_data[0]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[7]~0 (
	.dataa(src_data_151),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[7]~0_combout ),
	.cout());
defparam \av_ld_byte1_data[7]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[7]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[6]~1 (
	.dataa(src_data_14),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[6]~1_combout ),
	.cout());
defparam \av_ld_byte1_data[6]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[6]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[5]~2 (
	.dataa(src_data_131),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[5]~2_combout ),
	.cout());
defparam \av_ld_byte1_data[5]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[5]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[4]~3 (
	.dataa(src_data_121),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[4]~3_combout ),
	.cout());
defparam \av_ld_byte1_data[4]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[4]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[3]~4 (
	.dataa(src_data_111),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[3]~4_combout ),
	.cout());
defparam \av_ld_byte1_data[3]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[2]~5 (
	.dataa(src_data_10),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[2]~5_combout ),
	.cout());
defparam \av_ld_byte1_data[2]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[1]~6 (
	.dataa(src_data_9),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[1]~6_combout ),
	.cout());
defparam \av_ld_byte1_data[1]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[1]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[0]~7 (
	.dataa(src_data_8),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[0]~7_combout ),
	.cout());
defparam \av_ld_byte1_data[0]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[27]~27 (
	.dataa(\Add1~88_combout ),
	.datab(\E_logic_result[27]~29_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[27]~27_combout ),
	.cout());
defparam \W_alu_result[27]~27 .lut_mask = 16'hAACC;
defparam \W_alu_result[27]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[28]~28 (
	.dataa(\Add1~90_combout ),
	.datab(\E_logic_result[28]~28_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[28]~28_combout ),
	.cout());
defparam \W_alu_result[28]~28 .lut_mask = 16'hAACC;
defparam \W_alu_result[28]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[29]~29 (
	.dataa(\Add1~92_combout ),
	.datab(\E_logic_result[29]~27_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[29]~29_combout ),
	.cout());
defparam \W_alu_result[29]~29 .lut_mask = 16'hAACC;
defparam \W_alu_result[29]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[30]~30 (
	.dataa(\Add1~94_combout ),
	.datab(\E_logic_result[30]~26_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[30]~30_combout ),
	.cout());
defparam \W_alu_result[30]~30 .lut_mask = 16'hAACC;
defparam \W_alu_result[30]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[31]~31 (
	.dataa(\Add1~96_combout ),
	.datab(\E_logic_result[31]~25_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[31]~31_combout ),
	.cout());
defparam \W_alu_result[31]~31 .lut_mask = 16'hAACC;
defparam \W_alu_result[31]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld_signed~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~1_combout ),
	.cout());
defparam \D_ctrl_ld_signed~1 .lut_mask = 16'hEEEE;
defparam \D_ctrl_ld_signed~1 .sum_lutc_input = "datac";

dffeas R_wr_dst_reg(
	.clk(wire_pll7_clk_0),
	.d(\D_wr_dst_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_wr_dst_reg~q ),
	.prn(vcc));
defparam R_wr_dst_reg.is_wysiwyg = "true";
defparam R_wr_dst_reg.power_up = "low";

cycloneive_lcell_comb W_rf_wren(
	.dataa(r_sync_rst),
	.datab(\W_valid~q ),
	.datac(\R_wr_dst_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wren~combout ),
	.cout());
defparam W_rf_wren.lut_mask = 16'hFEFE;
defparam W_rf_wren.sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte0_data_nxt[0]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[0]~0 (
	.dataa(\R_ctrl_br_cmp~q ),
	.datab(\W_cmp_result~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~0_combout ),
	.cout());
defparam \W_rf_wr_data[0]~0 .lut_mask = 16'hEEEE;
defparam \W_rf_wr_data[0]~0 .sum_lutc_input = "datac";

dffeas \W_control_rd_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\E_control_rd_data[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[0]~q ),
	.prn(vcc));
defparam \W_control_rd_data[0] .is_wysiwyg = "true";
defparam \W_control_rd_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[0]~1 (
	.dataa(\W_control_rd_data[0]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\R_ctrl_rd_ctl_reg~q ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~1_combout ),
	.cout());
defparam \W_rf_wr_data[0]~1 .lut_mask = 16'hACFF;
defparam \W_rf_wr_data[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[0]~2 (
	.dataa(\av_ld_byte0_data[0]~q ),
	.datab(\W_rf_wr_data[0]~0_combout ),
	.datac(\W_rf_wr_data[0]~1_combout ),
	.datad(\R_ctrl_ld~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~2_combout ),
	.cout());
defparam \W_rf_wr_data[0]~2 .lut_mask = 16'hFAFC;
defparam \W_rf_wr_data[0]~2 .sum_lutc_input = "datac";

dffeas \R_dst_regnum[0] (
	.clk(wire_pll7_clk_0),
	.d(\D_dst_regnum[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[0]~q ),
	.prn(vcc));
defparam \R_dst_regnum[0] .is_wysiwyg = "true";
defparam \R_dst_regnum[0] .power_up = "low";

dffeas \R_dst_regnum[1] (
	.clk(wire_pll7_clk_0),
	.d(\D_dst_regnum[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[1]~q ),
	.prn(vcc));
defparam \R_dst_regnum[1] .is_wysiwyg = "true";
defparam \R_dst_regnum[1] .power_up = "low";

dffeas \R_dst_regnum[2] (
	.clk(wire_pll7_clk_0),
	.d(\D_dst_regnum[2]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[2]~q ),
	.prn(vcc));
defparam \R_dst_regnum[2] .is_wysiwyg = "true";
defparam \R_dst_regnum[2] .power_up = "low";

dffeas \R_dst_regnum[3] (
	.clk(wire_pll7_clk_0),
	.d(\D_dst_regnum[3]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[3]~q ),
	.prn(vcc));
defparam \R_dst_regnum[3] .is_wysiwyg = "true";
defparam \R_dst_regnum[3] .power_up = "low";

dffeas \R_dst_regnum[4] (
	.clk(wire_pll7_clk_0),
	.d(\D_dst_regnum[4]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[4]~q ),
	.prn(vcc));
defparam \R_dst_regnum[4] .is_wysiwyg = "true";
defparam \R_dst_regnum[4] .power_up = "low";

dffeas \av_ld_byte0_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte0_data_nxt[1]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[1] .power_up = "low";

dffeas \W_control_rd_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\E_control_rd_data[1]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[1]~q ),
	.prn(vcc));
defparam \W_control_rd_data[1] .is_wysiwyg = "true";
defparam \W_control_rd_data[1] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[1]~3 (
	.dataa(\W_control_rd_data[1]~q ),
	.datab(\W_alu_result[1]~q ),
	.datac(gnd),
	.datad(\R_ctrl_rd_ctl_reg~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[1]~3_combout ),
	.cout());
defparam \W_rf_wr_data[1]~3 .lut_mask = 16'hAACC;
defparam \W_rf_wr_data[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[1]~4 (
	.dataa(\av_ld_byte0_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_rf_wr_data[1]~3_combout ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[1]~4_combout ),
	.cout());
defparam \W_rf_wr_data[1]~4 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[1]~4 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte0_data_nxt[2]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[2] .power_up = "low";

dffeas \W_control_rd_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\E_control_rd_data[2]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[2]~q ),
	.prn(vcc));
defparam \W_control_rd_data[2] .is_wysiwyg = "true";
defparam \W_control_rd_data[2] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[2]~5 (
	.dataa(\W_control_rd_data[2]~q ),
	.datab(W_alu_result_2),
	.datac(gnd),
	.datad(\R_ctrl_rd_ctl_reg~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[2]~5_combout ),
	.cout());
defparam \W_rf_wr_data[2]~5 .lut_mask = 16'hAACC;
defparam \W_rf_wr_data[2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[2]~6 (
	.dataa(\av_ld_byte0_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_rf_wr_data[2]~5_combout ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[2]~6_combout ),
	.cout());
defparam \W_rf_wr_data[2]~6 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[2]~6 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte0_data_nxt[3]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[3] .power_up = "low";

dffeas \W_control_rd_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\E_control_rd_data[3]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[3]~q ),
	.prn(vcc));
defparam \W_control_rd_data[3] .is_wysiwyg = "true";
defparam \W_control_rd_data[3] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[3]~7 (
	.dataa(\W_control_rd_data[3]~q ),
	.datab(W_alu_result_3),
	.datac(gnd),
	.datad(\R_ctrl_rd_ctl_reg~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[3]~7_combout ),
	.cout());
defparam \W_rf_wr_data[3]~7 .lut_mask = 16'hAACC;
defparam \W_rf_wr_data[3]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[3]~8 (
	.dataa(\av_ld_byte0_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_rf_wr_data[3]~7_combout ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[3]~8_combout ),
	.cout());
defparam \W_rf_wr_data[3]~8 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[3]~8 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte0_data_nxt[4]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[4] .power_up = "low";

dffeas \W_control_rd_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\E_control_rd_data[4]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[4]~q ),
	.prn(vcc));
defparam \W_control_rd_data[4] .is_wysiwyg = "true";
defparam \W_control_rd_data[4] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[4]~9 (
	.dataa(\W_control_rd_data[4]~q ),
	.datab(W_alu_result_4),
	.datac(gnd),
	.datad(\R_ctrl_rd_ctl_reg~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[4]~9_combout ),
	.cout());
defparam \W_rf_wr_data[4]~9 .lut_mask = 16'hAACC;
defparam \W_rf_wr_data[4]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[4]~10 (
	.dataa(\av_ld_byte0_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_rf_wr_data[4]~9_combout ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[4]~10_combout ),
	.cout());
defparam \W_rf_wr_data[4]~10 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[4]~10 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte0_data_nxt[5]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[5] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[5]~11 (
	.dataa(\av_ld_byte0_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_5),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[5]~11_combout ),
	.cout());
defparam \W_rf_wr_data[5]~11 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[5]~11 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte0_data_nxt[6]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[6] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[6]~12 (
	.dataa(\av_ld_byte0_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_6),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[6]~12_combout ),
	.cout());
defparam \W_rf_wr_data[6]~12 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[6]~12 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte0_data_nxt[7]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[7] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[7]~13 (
	.dataa(\av_ld_byte0_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_7),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[7]~13_combout ),
	.cout());
defparam \W_rf_wr_data[7]~13 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[7]~13 .sum_lutc_input = "datac";

dffeas \D_iw[31] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[31]~77_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

dffeas \av_ld_byte3_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte3_data_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[2] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[26]~14 (
	.dataa(\av_ld_byte3_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_26),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[26]~14_combout ),
	.cout());
defparam \W_rf_wr_data[26]~14 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[26]~14 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte3_data_nxt~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[1] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[25]~15 (
	.dataa(\av_ld_byte3_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_25),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[25]~15_combout ),
	.cout());
defparam \W_rf_wr_data[25]~15 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[25]~15 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte3_data_nxt~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[24]~16 (
	.dataa(\av_ld_byte3_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_24),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[24]~16_combout ),
	.cout());
defparam \W_rf_wr_data[24]~16 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[24]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[23]~17 (
	.dataa(\av_ld_byte2_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_23),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[23]~17_combout ),
	.cout());
defparam \W_rf_wr_data[23]~17 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[23]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[22]~18 (
	.dataa(\av_ld_byte2_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_22),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[22]~18_combout ),
	.cout());
defparam \W_rf_wr_data[22]~18 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[22]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[21]~19 (
	.dataa(\av_ld_byte2_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_21),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[21]~19_combout ),
	.cout());
defparam \W_rf_wr_data[21]~19 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[21]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[20]~20 (
	.dataa(\av_ld_byte2_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_20),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[20]~20_combout ),
	.cout());
defparam \W_rf_wr_data[20]~20 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[20]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[19]~21 (
	.dataa(\av_ld_byte2_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_19),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[19]~21_combout ),
	.cout());
defparam \W_rf_wr_data[19]~21 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[19]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[18]~22 (
	.dataa(\av_ld_byte2_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_18),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[18]~22_combout ),
	.cout());
defparam \W_rf_wr_data[18]~22 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[18]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[17]~23 (
	.dataa(\av_ld_byte2_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_17),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[17]~23_combout ),
	.cout());
defparam \W_rf_wr_data[17]~23 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[17]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[16]~24 (
	.dataa(\av_ld_byte2_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_16),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[16]~24_combout ),
	.cout());
defparam \W_rf_wr_data[16]~24 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[16]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[15]~25 (
	.dataa(\av_ld_byte1_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_15),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[15]~25_combout ),
	.cout());
defparam \W_rf_wr_data[15]~25 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[15]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[14]~26 (
	.dataa(\av_ld_byte1_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_14),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[14]~26_combout ),
	.cout());
defparam \W_rf_wr_data[14]~26 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[14]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[13]~27 (
	.dataa(\av_ld_byte1_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_13),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[13]~27_combout ),
	.cout());
defparam \W_rf_wr_data[13]~27 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[13]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[12]~28 (
	.dataa(\av_ld_byte1_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_12),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[12]~28_combout ),
	.cout());
defparam \W_rf_wr_data[12]~28 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[12]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[11]~29 (
	.dataa(\av_ld_byte1_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_11),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[11]~29_combout ),
	.cout());
defparam \W_rf_wr_data[11]~29 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[11]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[10]~30 (
	.dataa(\av_ld_byte1_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_10),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[10]~30_combout ),
	.cout());
defparam \W_rf_wr_data[10]~30 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[10]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[9]~31 (
	.dataa(\av_ld_byte1_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_9),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[9]~31_combout ),
	.cout());
defparam \W_rf_wr_data[9]~31 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[9]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[8]~32 (
	.dataa(\av_ld_byte1_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_8),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[8]~32_combout ),
	.cout());
defparam \W_rf_wr_data[8]~32 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[8]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~0 (
	.dataa(\Equal0~16_combout ),
	.datab(\Equal0~14_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~0_combout ),
	.cout());
defparam \D_wr_dst_reg~0 .lut_mask = 16'hEFFF;
defparam \D_wr_dst_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~1 (
	.dataa(\Equal0~17_combout ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\R_ctrl_br_nxt~0_combout ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~1_combout ),
	.cout());
defparam \D_wr_dst_reg~1 .lut_mask = 16'hFEFF;
defparam \D_wr_dst_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[1]~0 (
	.dataa(\D_iw[23]~q ),
	.datab(\D_iw[18]~q ),
	.datac(gnd),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~0_combout ),
	.cout());
defparam \D_dst_regnum[1]~0 .lut_mask = 16'hAACC;
defparam \D_dst_regnum[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~3 (
	.dataa(\Equal62~10_combout ),
	.datab(\Equal62~13_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~3 .lut_mask = 16'hEFFE;
defparam \D_ctrl_implicit_dst_eretaddr~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~4 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~4 .lut_mask = 16'hFBFF;
defparam \D_ctrl_implicit_dst_eretaddr~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~5 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datac(\D_ctrl_exception~11_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~5 .lut_mask = 16'hFFFE;
defparam \D_ctrl_implicit_dst_eretaddr~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~6 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.datab(\D_ctrl_exception~17_combout ),
	.datac(\D_ctrl_exception~21_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~6_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~6 .lut_mask = 16'hBFFF;
defparam \D_ctrl_implicit_dst_eretaddr~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[1]~1 (
	.dataa(\Equal0~4_combout ),
	.datab(\D_ctrl_jmp_direct~0_combout ),
	.datac(\D_dst_regnum[1]~0_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~6_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~1_combout ),
	.cout());
defparam \D_dst_regnum[1]~1 .lut_mask = 16'hFEFF;
defparam \D_dst_regnum[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[2]~2 (
	.dataa(\Equal0~14_combout ),
	.datab(\D_iw[4]~q ),
	.datac(\Equal0~4_combout ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[2]~2_combout ),
	.cout());
defparam \D_dst_regnum[2]~2 .lut_mask = 16'hDF1F;
defparam \D_dst_regnum[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[2]~3 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.datab(\D_ctrl_force_src2_zero~0_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_dst_regnum[2]~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[2]~3_combout ),
	.cout());
defparam \D_dst_regnum[2]~3 .lut_mask = 16'hFFDF;
defparam \D_dst_regnum[2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[2]~4 (
	.dataa(\D_ctrl_exception~17_combout ),
	.datab(\D_ctrl_exception~21_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datad(\D_dst_regnum[2]~3_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[2]~4_combout ),
	.cout());
defparam \D_dst_regnum[2]~4 .lut_mask = 16'hFFFE;
defparam \D_dst_regnum[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[2]~5 (
	.dataa(\D_iw[24]~q ),
	.datab(\D_iw[19]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\D_dst_regnum[2]~4_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[2]~5_combout ),
	.cout());
defparam \D_dst_regnum[2]~5 .lut_mask = 16'hACFF;
defparam \D_dst_regnum[2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~6 (
	.dataa(\D_iw[26]~q ),
	.datab(\D_iw[21]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\D_dst_regnum[2]~4_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~6_combout ),
	.cout());
defparam \D_dst_regnum[4]~6 .lut_mask = 16'hACFF;
defparam \D_dst_regnum[4]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[3]~7 (
	.dataa(\D_iw[25]~q ),
	.datab(\D_iw[20]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\D_dst_regnum[2]~4_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[3]~7_combout ),
	.cout());
defparam \D_dst_regnum[3]~7 .lut_mask = 16'hACFF;
defparam \D_dst_regnum[3]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~19 (
	.dataa(\D_dst_regnum[1]~1_combout ),
	.datab(\D_dst_regnum[2]~5_combout ),
	.datac(\D_dst_regnum[4]~6_combout ),
	.datad(\D_dst_regnum[3]~7_combout ),
	.cin(gnd),
	.combout(\Equal0~19_combout ),
	.cout());
defparam \Equal0~19 .lut_mask = 16'h7FFF;
defparam \Equal0~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~8 (
	.dataa(\D_iw[22]~q ),
	.datab(\D_iw[17]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\D_dst_regnum[2]~4_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~8_combout ),
	.cout());
defparam \D_dst_regnum[0]~8 .lut_mask = 16'hACFF;
defparam \D_dst_regnum[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~2 (
	.dataa(\D_wr_dst_reg~0_combout ),
	.datab(\D_wr_dst_reg~1_combout ),
	.datac(\Equal0~19_combout ),
	.datad(\D_dst_regnum[0]~8_combout ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~2_combout ),
	.cout());
defparam \D_wr_dst_reg~2 .lut_mask = 16'hFF7F;
defparam \D_wr_dst_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_rshift8~0 (
	.dataa(\W_alu_result[1]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\av_ld_align_cycle[0]~q ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_rshift8~0_combout ),
	.cout());
defparam \av_ld_rshift8~0 .lut_mask = 16'hEFFF;
defparam \av_ld_rshift8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_rshift8~1 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_rshift8~1_combout ),
	.cout());
defparam \av_ld_rshift8~1 .lut_mask = 16'hEEEE;
defparam \av_ld_rshift8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data[2]~0 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\av_ld_rshift8~0_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data[2]~0_combout ),
	.cout());
defparam \av_ld_byte0_data[2]~0 .lut_mask = 16'hFF55;
defparam \av_ld_byte0_data[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~0 (
	.dataa(\E_wrctl_status~0_combout ),
	.datab(\W_ipending_reg[0]~q ),
	.datac(\W_status_reg_pie~q ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~0_combout ),
	.cout());
defparam \E_control_rd_data[0]~0 .lut_mask = 16'hFAFC;
defparam \E_control_rd_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~1 (
	.dataa(\W_estatus_reg~q ),
	.datab(\W_bstatus_reg~q ),
	.datac(\D_iw[7]~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~1_combout ),
	.cout());
defparam \E_control_rd_data[0]~1 .lut_mask = 16'hEFFE;
defparam \E_control_rd_data[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~2 (
	.dataa(\Equal135~0_combout ),
	.datab(\E_control_rd_data[0]~0_combout ),
	.datac(\E_control_rd_data[0]~1_combout ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~2_combout ),
	.cout());
defparam \E_control_rd_data[0]~2 .lut_mask = 16'hFEFF;
defparam \E_control_rd_data[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~3 (
	.dataa(\E_control_rd_data[0]~2_combout ),
	.datab(\W_ienable_reg[0]~q ),
	.datac(\Equal135~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~3_combout ),
	.cout());
defparam \E_control_rd_data[0]~3 .lut_mask = 16'hFEFE;
defparam \E_control_rd_data[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_control_rd_data[1]~0 (
	.dataa(\D_iw[8]~q ),
	.datab(\D_iw[7]~q ),
	.datac(\D_iw[6]~q ),
	.datad(\Equal135~0_combout ),
	.cin(gnd),
	.combout(\W_control_rd_data[1]~0_combout ),
	.cout());
defparam \W_control_rd_data[1]~0 .lut_mask = 16'h96FF;
defparam \W_control_rd_data[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[1]~4 (
	.dataa(\W_ienable_reg[1]~q ),
	.datab(\W_ipending_reg[1]~q ),
	.datac(\Equal135~1_combout ),
	.datad(\W_control_rd_data[1]~0_combout ),
	.cin(gnd),
	.combout(\E_control_rd_data[1]~4_combout ),
	.cout());
defparam \E_control_rd_data[1]~4 .lut_mask = 16'hACFF;
defparam \E_control_rd_data[1]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[2]~14 (
	.dataa(\av_ld_byte1_data[2]~q ),
	.datab(src_data_2),
	.datac(src_data_21),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~14_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~14 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[2]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[2]~5 (
	.dataa(\W_ienable_reg[2]~q ),
	.datab(\W_ipending_reg[2]~q ),
	.datac(\Equal135~1_combout ),
	.datad(\W_control_rd_data[1]~0_combout ),
	.cin(gnd),
	.combout(\E_control_rd_data[2]~5_combout ),
	.cout());
defparam \E_control_rd_data[2]~5 .lut_mask = 16'hACFF;
defparam \E_control_rd_data[2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[3]~6 (
	.dataa(\W_ienable_reg[3]~q ),
	.datab(\W_ipending_reg[3]~q ),
	.datac(\Equal135~1_combout ),
	.datad(\W_control_rd_data[1]~0_combout ),
	.cin(gnd),
	.combout(\E_control_rd_data[3]~6_combout ),
	.cout());
defparam \E_control_rd_data[3]~6 .lut_mask = 16'hACFF;
defparam \E_control_rd_data[3]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[4]~7 (
	.dataa(\W_ienable_reg[4]~q ),
	.datab(\W_ipending_reg[4]~q ),
	.datac(\Equal135~1_combout ),
	.datad(\W_control_rd_data[1]~0_combout ),
	.cin(gnd),
	.combout(\E_control_rd_data[4]~7_combout ),
	.cout());
defparam \E_control_rd_data[4]~7 .lut_mask = 16'hACFF;
defparam \E_control_rd_data[4]~7 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte3_data_nxt~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[3] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[27]~33 (
	.dataa(\av_ld_byte3_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[27]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[27]~33_combout ),
	.cout());
defparam \W_rf_wr_data[27]~33 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[27]~33 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte3_data_nxt~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[4] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[28]~34 (
	.dataa(\av_ld_byte3_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[28]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[28]~34_combout ),
	.cout());
defparam \W_rf_wr_data[28]~34 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[28]~34 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte3_data_nxt~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[5] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[29]~35 (
	.dataa(\av_ld_byte3_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[29]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[29]~35_combout ),
	.cout());
defparam \W_rf_wr_data[29]~35 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[29]~35 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte3_data_nxt~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[6] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[30]~36 (
	.dataa(\av_ld_byte3_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[30]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[30]~36_combout ),
	.cout());
defparam \W_rf_wr_data[30]~36 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[30]~36 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_byte3_data_nxt~35_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[7] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[31]~37 (
	.dataa(\av_ld_byte3_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[31]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[31]~37_combout ),
	.cout());
defparam \W_rf_wr_data[31]~37 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[31]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[31]~76 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_31),
	.datad(out_data_buffer_31),
	.cin(gnd),
	.combout(\F_iw[31]~76_combout ),
	.cout());
defparam \F_iw[31]~76 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[31]~77 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[31]~76_combout ),
	.datac(src_payload),
	.datad(out_payload_15),
	.cin(gnd),
	.combout(\F_iw[31]~77_combout ),
	.cout());
defparam \F_iw[31]~77 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~77 .sum_lutc_input = "datac";

dffeas R_ctrl_ld_signed(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_ld_signed~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld_signed~q ),
	.prn(vcc));
defparam R_ctrl_ld_signed.is_wysiwyg = "true";
defparam R_ctrl_ld_signed.power_up = "low";

cycloneive_lcell_comb \av_fill_bit~0 (
	.dataa(\R_ctrl_ld_signed~q ),
	.datab(\av_ld_byte1_data[7]~q ),
	.datac(\av_ld_byte0_data[7]~q ),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\av_fill_bit~0_combout ),
	.cout());
defparam \av_fill_bit~0 .lut_mask = 16'hFAFC;
defparam \av_fill_bit~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~0 (
	.dataa(source_addr_1),
	.datab(src0_valid),
	.datac(out_payload_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~0_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~0 .lut_mask = 16'hFEFE;
defparam \av_ld_byte3_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~1 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_26),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~1_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~1 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~2 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_01),
	.datac(readdata_26),
	.datad(av_readdata_pre_301),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~2_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~2 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~3 (
	.dataa(\av_ld_byte3_data_nxt~1_combout ),
	.datab(\av_ld_byte3_data_nxt~2_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_261),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~3_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~3 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~4 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~0_combout ),
	.datac(\av_ld_byte3_data_nxt~3_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~4_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~4 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~5 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_25),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~5_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~5 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~6 (
	.dataa(out_valid1),
	.datab(read_latency_shift_reg_01),
	.datac(readdata_25),
	.datad(out_data_buffer_251),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~6_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~6 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~7 (
	.dataa(\av_ld_byte3_data_nxt~5_combout ),
	.datab(\av_ld_byte3_data_nxt~6_combout ),
	.datac(out_payload_9),
	.datad(src_payload3),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~7_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~7 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~8 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~7_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~8_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~8 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~9 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_24),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~9_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~9 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~10 (
	.dataa(out_valid1),
	.datab(read_latency_shift_reg_01),
	.datac(readdata_24),
	.datad(out_data_buffer_241),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~10_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~10 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~11 (
	.dataa(\av_ld_byte3_data_nxt~9_combout ),
	.datab(\av_ld_byte3_data_nxt~10_combout ),
	.datac(out_payload_8),
	.datad(src_payload3),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~11_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~11 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~12 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~11_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~12_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~12 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data_en~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\D_ctrl_mem16~0_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data_en~0_combout ),
	.cout());
defparam \av_ld_byte1_data_en~0 .lut_mask = 16'hEFFF;
defparam \av_ld_byte1_data_en~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~13 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_27),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~13_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~13 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~14 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_01),
	.datac(readdata_271),
	.datad(av_readdata_pre_301),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~14_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~14 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~15 (
	.dataa(\av_ld_byte3_data_nxt~13_combout ),
	.datab(\av_ld_byte3_data_nxt~14_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_271),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~15_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~15 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~16 (
	.dataa(\av_ld_byte3_data_nxt~15_combout ),
	.datab(source_addr_1),
	.datac(src0_valid),
	.datad(out_payload_11),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~16_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~16 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~17 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~16_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~17_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~17 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~18 (
	.dataa(source_addr_1),
	.datab(src0_valid),
	.datac(out_payload_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~18_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~18 .lut_mask = 16'hFEFE;
defparam \av_ld_byte3_data_nxt~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~19 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_28),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~19_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~19 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~20 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_01),
	.datac(readdata_281),
	.datad(av_readdata_pre_301),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~20_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~20 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~21 (
	.dataa(\av_ld_byte3_data_nxt~19_combout ),
	.datab(\av_ld_byte3_data_nxt~20_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_281),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~21_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~21 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~22 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~18_combout ),
	.datac(\av_ld_byte3_data_nxt~21_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~22_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~22 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~23 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_29),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~23_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~23 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~24 (
	.dataa(out_valid1),
	.datab(read_latency_shift_reg_01),
	.datac(readdata_291),
	.datad(out_data_buffer_291),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~24_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~24 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~25 (
	.dataa(\av_ld_byte3_data_nxt~23_combout ),
	.datab(\av_ld_byte3_data_nxt~24_combout ),
	.datac(out_payload_13),
	.datad(src_payload3),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~25_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~25 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~26 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~25_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~26_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~26 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~27 (
	.dataa(source_addr_1),
	.datab(src0_valid),
	.datac(out_payload_14),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~27_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~27 .lut_mask = 16'hFEFE;
defparam \av_ld_byte3_data_nxt~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~28 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_30),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~28_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~28 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~29 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_01),
	.datac(readdata_301),
	.datad(av_readdata_pre_301),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~29_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~29 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~30 (
	.dataa(\av_ld_byte3_data_nxt~28_combout ),
	.datab(\av_ld_byte3_data_nxt~29_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_301),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~30_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~30 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~31 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~27_combout ),
	.datac(\av_ld_byte3_data_nxt~30_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~31_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~31 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~32 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_31),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~32_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~32 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~33 (
	.dataa(out_valid1),
	.datab(read_latency_shift_reg_01),
	.datac(readdata_31),
	.datad(out_data_buffer_311),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~33_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~33 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~34 (
	.dataa(\av_ld_byte3_data_nxt~32_combout ),
	.datab(\av_ld_byte3_data_nxt~33_combout ),
	.datac(out_payload_15),
	.datad(src_payload3),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~34_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~34 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~35 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~34_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~35_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~35 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[0]~15 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[0]~q ),
	.datad(src_data_0),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[0]~15_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[0]~15 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[0]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[1]~16 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[1]~q ),
	.datad(src_data_12),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~16_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~16 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[1]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[3]~17 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[3]~q ),
	.datad(src_data_31),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~17_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~17 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[3]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[4]~18 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[4]~q ),
	.datad(src_data_41),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~18_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~18 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[4]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[5]~19 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[5]~q ),
	.datad(src_data_51),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~19_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~19 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[5]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[6]~20 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[6]~q ),
	.datad(src_data_6),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~20_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~20 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[6]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[7]~21 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[7]~q ),
	.datad(src_data_7),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~21_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~21 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[7]~21 .sum_lutc_input = "datac";

dffeas \W_alu_result[6] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[6]~20_combout ),
	.asdata(\E_shift_rot_result[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_6),
	.prn(vcc));
defparam \W_alu_result[6] .is_wysiwyg = "true";
defparam \W_alu_result[6] .power_up = "low";

dffeas \W_alu_result[26] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[26]~0_combout ),
	.asdata(\E_shift_rot_result[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_26),
	.prn(vcc));
defparam \W_alu_result[26] .is_wysiwyg = "true";
defparam \W_alu_result[26] .power_up = "low";

dffeas \W_alu_result[25] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[25]~1_combout ),
	.asdata(\E_shift_rot_result[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_25),
	.prn(vcc));
defparam \W_alu_result[25] .is_wysiwyg = "true";
defparam \W_alu_result[25] .power_up = "low";

dffeas \W_alu_result[24] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[24]~2_combout ),
	.asdata(\E_shift_rot_result[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_24),
	.prn(vcc));
defparam \W_alu_result[24] .is_wysiwyg = "true";
defparam \W_alu_result[24] .power_up = "low";

dffeas \W_alu_result[23] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[23]~3_combout ),
	.asdata(\E_shift_rot_result[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_23),
	.prn(vcc));
defparam \W_alu_result[23] .is_wysiwyg = "true";
defparam \W_alu_result[23] .power_up = "low";

dffeas \W_alu_result[22] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[22]~4_combout ),
	.asdata(\E_shift_rot_result[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_22),
	.prn(vcc));
defparam \W_alu_result[22] .is_wysiwyg = "true";
defparam \W_alu_result[22] .power_up = "low";

dffeas \W_alu_result[21] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[21]~5_combout ),
	.asdata(\E_shift_rot_result[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_21),
	.prn(vcc));
defparam \W_alu_result[21] .is_wysiwyg = "true";
defparam \W_alu_result[21] .power_up = "low";

dffeas \W_alu_result[20] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[20]~6_combout ),
	.asdata(\E_shift_rot_result[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_20),
	.prn(vcc));
defparam \W_alu_result[20] .is_wysiwyg = "true";
defparam \W_alu_result[20] .power_up = "low";

dffeas \W_alu_result[19] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[19]~7_combout ),
	.asdata(\E_shift_rot_result[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_19),
	.prn(vcc));
defparam \W_alu_result[19] .is_wysiwyg = "true";
defparam \W_alu_result[19] .power_up = "low";

dffeas \W_alu_result[18] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[18]~8_combout ),
	.asdata(\E_shift_rot_result[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_18),
	.prn(vcc));
defparam \W_alu_result[18] .is_wysiwyg = "true";
defparam \W_alu_result[18] .power_up = "low";

dffeas \W_alu_result[17] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[17]~9_combout ),
	.asdata(\E_shift_rot_result[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_17),
	.prn(vcc));
defparam \W_alu_result[17] .is_wysiwyg = "true";
defparam \W_alu_result[17] .power_up = "low";

dffeas \W_alu_result[16] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[16]~10_combout ),
	.asdata(\E_shift_rot_result[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_16),
	.prn(vcc));
defparam \W_alu_result[16] .is_wysiwyg = "true";
defparam \W_alu_result[16] .power_up = "low";

dffeas \W_alu_result[15] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[15]~11_combout ),
	.asdata(\E_shift_rot_result[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_15),
	.prn(vcc));
defparam \W_alu_result[15] .is_wysiwyg = "true";
defparam \W_alu_result[15] .power_up = "low";

dffeas \W_alu_result[14] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[14]~12_combout ),
	.asdata(\E_shift_rot_result[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_14),
	.prn(vcc));
defparam \W_alu_result[14] .is_wysiwyg = "true";
defparam \W_alu_result[14] .power_up = "low";

dffeas \W_alu_result[13] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[13]~13_combout ),
	.asdata(\E_shift_rot_result[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_13),
	.prn(vcc));
defparam \W_alu_result[13] .is_wysiwyg = "true";
defparam \W_alu_result[13] .power_up = "low";

dffeas \W_alu_result[12] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[12]~14_combout ),
	.asdata(\E_shift_rot_result[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_12),
	.prn(vcc));
defparam \W_alu_result[12] .is_wysiwyg = "true";
defparam \W_alu_result[12] .power_up = "low";

dffeas \W_alu_result[11] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[11]~15_combout ),
	.asdata(\E_shift_rot_result[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_11),
	.prn(vcc));
defparam \W_alu_result[11] .is_wysiwyg = "true";
defparam \W_alu_result[11] .power_up = "low";

dffeas \W_alu_result[10] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[10]~16_combout ),
	.asdata(\E_shift_rot_result[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_10),
	.prn(vcc));
defparam \W_alu_result[10] .is_wysiwyg = "true";
defparam \W_alu_result[10] .power_up = "low";

dffeas \W_alu_result[5] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[5]~21_combout ),
	.asdata(\E_shift_rot_result[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_5),
	.prn(vcc));
defparam \W_alu_result[5] .is_wysiwyg = "true";
defparam \W_alu_result[5] .power_up = "low";

dffeas \W_alu_result[7] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[7]~19_combout ),
	.asdata(\E_shift_rot_result[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_7),
	.prn(vcc));
defparam \W_alu_result[7] .is_wysiwyg = "true";
defparam \W_alu_result[7] .power_up = "low";

dffeas \W_alu_result[9] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[9]~17_combout ),
	.asdata(\E_shift_rot_result[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_9),
	.prn(vcc));
defparam \W_alu_result[9] .is_wysiwyg = "true";
defparam \W_alu_result[9] .power_up = "low";

dffeas \W_alu_result[8] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[8]~18_combout ),
	.asdata(\E_shift_rot_result[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_8),
	.prn(vcc));
defparam \W_alu_result[8] .is_wysiwyg = "true";
defparam \W_alu_result[8] .power_up = "low";

dffeas \W_alu_result[4] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[4]~22_combout ),
	.asdata(\E_shift_rot_result[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_4),
	.prn(vcc));
defparam \W_alu_result[4] .is_wysiwyg = "true";
defparam \W_alu_result[4] .power_up = "low";

dffeas \W_alu_result[3] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[3]~23_combout ),
	.asdata(\E_shift_rot_result[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_3),
	.prn(vcc));
defparam \W_alu_result[3] .is_wysiwyg = "true";
defparam \W_alu_result[3] .power_up = "low";

dffeas \W_alu_result[2] (
	.clk(wire_pll7_clk_0),
	.d(\W_alu_result[2]~24_combout ),
	.asdata(\E_shift_rot_result[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_2),
	.prn(vcc));
defparam \W_alu_result[2] .is_wysiwyg = "true";
defparam \W_alu_result[2] .power_up = "low";

dffeas \d_writedata[24] (
	.clk(wire_pll7_clk_0),
	.d(\d_writedata[24]~0_combout ),
	.asdata(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_24),
	.prn(vcc));
defparam \d_writedata[24] .is_wysiwyg = "true";
defparam \d_writedata[24] .power_up = "low";

dffeas \d_writedata[25] (
	.clk(wire_pll7_clk_0),
	.d(\d_writedata[25]~1_combout ),
	.asdata(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_25),
	.prn(vcc));
defparam \d_writedata[25] .is_wysiwyg = "true";
defparam \d_writedata[25] .power_up = "low";

dffeas \d_writedata[26] (
	.clk(wire_pll7_clk_0),
	.d(\d_writedata[26]~2_combout ),
	.asdata(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_26),
	.prn(vcc));
defparam \d_writedata[26] .is_wysiwyg = "true";
defparam \d_writedata[26] .power_up = "low";

dffeas \d_writedata[27] (
	.clk(wire_pll7_clk_0),
	.d(\d_writedata[27]~3_combout ),
	.asdata(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_27),
	.prn(vcc));
defparam \d_writedata[27] .is_wysiwyg = "true";
defparam \d_writedata[27] .power_up = "low";

dffeas \d_writedata[28] (
	.clk(wire_pll7_clk_0),
	.d(\d_writedata[28]~4_combout ),
	.asdata(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_28),
	.prn(vcc));
defparam \d_writedata[28] .is_wysiwyg = "true";
defparam \d_writedata[28] .power_up = "low";

dffeas \d_writedata[29] (
	.clk(wire_pll7_clk_0),
	.d(\d_writedata[29]~5_combout ),
	.asdata(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_29),
	.prn(vcc));
defparam \d_writedata[29] .is_wysiwyg = "true";
defparam \d_writedata[29] .power_up = "low";

dffeas \d_writedata[30] (
	.clk(wire_pll7_clk_0),
	.d(\d_writedata[30]~6_combout ),
	.asdata(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_30),
	.prn(vcc));
defparam \d_writedata[30] .is_wysiwyg = "true";
defparam \d_writedata[30] .power_up = "low";

dffeas \d_writedata[31] (
	.clk(wire_pll7_clk_0),
	.d(\d_writedata[31]~7_combout ),
	.asdata(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_31),
	.prn(vcc));
defparam \d_writedata[31] .is_wysiwyg = "true";
defparam \d_writedata[31] .power_up = "low";

dffeas d_read(
	.clk(wire_pll7_clk_0),
	.d(\d_read_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

dffeas d_write(
	.clk(wire_pll7_clk_0),
	.d(\E_st_stall~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas \d_writedata[0] (
	.clk(wire_pll7_clk_0),
	.d(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_0),
	.prn(vcc));
defparam \d_writedata[0] .is_wysiwyg = "true";
defparam \d_writedata[0] .power_up = "low";

dffeas \d_byteenable[0] (
	.clk(wire_pll7_clk_0),
	.d(\E_mem_byte_en[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_0),
	.prn(vcc));
defparam \d_byteenable[0] .is_wysiwyg = "true";
defparam \d_byteenable[0] .power_up = "low";

dffeas \d_writedata[1] (
	.clk(wire_pll7_clk_0),
	.d(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_1),
	.prn(vcc));
defparam \d_writedata[1] .is_wysiwyg = "true";
defparam \d_writedata[1] .power_up = "low";

dffeas \d_writedata[2] (
	.clk(wire_pll7_clk_0),
	.d(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_2),
	.prn(vcc));
defparam \d_writedata[2] .is_wysiwyg = "true";
defparam \d_writedata[2] .power_up = "low";

dffeas \d_writedata[3] (
	.clk(wire_pll7_clk_0),
	.d(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_3),
	.prn(vcc));
defparam \d_writedata[3] .is_wysiwyg = "true";
defparam \d_writedata[3] .power_up = "low";

dffeas \d_writedata[4] (
	.clk(wire_pll7_clk_0),
	.d(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_4),
	.prn(vcc));
defparam \d_writedata[4] .is_wysiwyg = "true";
defparam \d_writedata[4] .power_up = "low";

dffeas \d_writedata[5] (
	.clk(wire_pll7_clk_0),
	.d(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_5),
	.prn(vcc));
defparam \d_writedata[5] .is_wysiwyg = "true";
defparam \d_writedata[5] .power_up = "low";

dffeas \d_writedata[6] (
	.clk(wire_pll7_clk_0),
	.d(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_6),
	.prn(vcc));
defparam \d_writedata[6] .is_wysiwyg = "true";
defparam \d_writedata[6] .power_up = "low";

dffeas \d_writedata[7] (
	.clk(wire_pll7_clk_0),
	.d(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_7),
	.prn(vcc));
defparam \d_writedata[7] .is_wysiwyg = "true";
defparam \d_writedata[7] .power_up = "low";

dffeas \d_byteenable[1] (
	.clk(wire_pll7_clk_0),
	.d(\E_mem_byte_en[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_1),
	.prn(vcc));
defparam \d_byteenable[1] .is_wysiwyg = "true";
defparam \d_byteenable[1] .power_up = "low";

dffeas i_read(
	.clk(wire_pll7_clk_0),
	.d(\i_read_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas \F_pc[24] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[24]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_24),
	.prn(vcc));
defparam \F_pc[24] .is_wysiwyg = "true";
defparam \F_pc[24] .power_up = "low";

dffeas \F_pc[23] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[23]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_23),
	.prn(vcc));
defparam \F_pc[23] .is_wysiwyg = "true";
defparam \F_pc[23] .power_up = "low";

dffeas \F_pc[22] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[22]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_22),
	.prn(vcc));
defparam \F_pc[22] .is_wysiwyg = "true";
defparam \F_pc[22] .power_up = "low";

dffeas \F_pc[21] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[21]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_21),
	.prn(vcc));
defparam \F_pc[21] .is_wysiwyg = "true";
defparam \F_pc[21] .power_up = "low";

dffeas \F_pc[20] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[20]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_20),
	.prn(vcc));
defparam \F_pc[20] .is_wysiwyg = "true";
defparam \F_pc[20] .power_up = "low";

dffeas \F_pc[19] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[19]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_19),
	.prn(vcc));
defparam \F_pc[19] .is_wysiwyg = "true";
defparam \F_pc[19] .power_up = "low";

dffeas \F_pc[18] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[18]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_18),
	.prn(vcc));
defparam \F_pc[18] .is_wysiwyg = "true";
defparam \F_pc[18] .power_up = "low";

dffeas \F_pc[17] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[17]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_17),
	.prn(vcc));
defparam \F_pc[17] .is_wysiwyg = "true";
defparam \F_pc[17] .power_up = "low";

dffeas \F_pc[16] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[16]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_16),
	.prn(vcc));
defparam \F_pc[16] .is_wysiwyg = "true";
defparam \F_pc[16] .power_up = "low";

dffeas \F_pc[15] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[15]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_15),
	.prn(vcc));
defparam \F_pc[15] .is_wysiwyg = "true";
defparam \F_pc[15] .power_up = "low";

dffeas \F_pc[14] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[14]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_14),
	.prn(vcc));
defparam \F_pc[14] .is_wysiwyg = "true";
defparam \F_pc[14] .power_up = "low";

dffeas \F_pc[13] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[13]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_13),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

dffeas \F_pc[12] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[12]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_12),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

dffeas \F_pc[11] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[11]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_11),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

dffeas \F_pc[10] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[10]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_10),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

dffeas \F_pc[8] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[8]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_8),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

dffeas \F_pc[9] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[9]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_9),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

dffeas \F_pc[0] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[0]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_0),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

dffeas \F_pc[1] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[1]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_1),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

dffeas \F_pc[2] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[2]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_2),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

dffeas \F_pc[3] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[3]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_3),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

dffeas \F_pc[4] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[4]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_4),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

dffeas \F_pc[5] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[5]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_5),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

dffeas \F_pc[6] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[6]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_6),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

dffeas \F_pc[7] (
	.clk(wire_pll7_clk_0),
	.d(\F_pc_no_crst_nxt[7]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_7),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

dffeas \d_writedata[10] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[10]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_10),
	.prn(vcc));
defparam \d_writedata[10] .is_wysiwyg = "true";
defparam \d_writedata[10] .power_up = "low";

dffeas \d_byteenable[2] (
	.clk(wire_pll7_clk_0),
	.d(\E_mem_byte_en[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_2),
	.prn(vcc));
defparam \d_byteenable[2] .is_wysiwyg = "true";
defparam \d_byteenable[2] .power_up = "low";

dffeas \d_byteenable[3] (
	.clk(wire_pll7_clk_0),
	.d(\E_mem_byte_en[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_3),
	.prn(vcc));
defparam \d_byteenable[3] .is_wysiwyg = "true";
defparam \d_byteenable[3] .power_up = "low";

dffeas hbreak_enabled(
	.clk(wire_pll7_clk_0),
	.d(\hbreak_enabled~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas \d_writedata[8] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[8]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_8),
	.prn(vcc));
defparam \d_writedata[8] .is_wysiwyg = "true";
defparam \d_writedata[8] .power_up = "low";

dffeas \d_writedata[9] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[9]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_9),
	.prn(vcc));
defparam \d_writedata[9] .is_wysiwyg = "true";
defparam \d_writedata[9] .power_up = "low";

dffeas \d_writedata[11] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[11]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_11),
	.prn(vcc));
defparam \d_writedata[11] .is_wysiwyg = "true";
defparam \d_writedata[11] .power_up = "low";

dffeas \d_writedata[12] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[12]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_12),
	.prn(vcc));
defparam \d_writedata[12] .is_wysiwyg = "true";
defparam \d_writedata[12] .power_up = "low";

dffeas \d_writedata[13] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[13]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_13),
	.prn(vcc));
defparam \d_writedata[13] .is_wysiwyg = "true";
defparam \d_writedata[13] .power_up = "low";

dffeas \d_writedata[14] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[14]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_14),
	.prn(vcc));
defparam \d_writedata[14] .is_wysiwyg = "true";
defparam \d_writedata[14] .power_up = "low";

dffeas \d_writedata[15] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[15]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_15),
	.prn(vcc));
defparam \d_writedata[15] .is_wysiwyg = "true";
defparam \d_writedata[15] .power_up = "low";

dffeas \d_writedata[16] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[16]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_16),
	.prn(vcc));
defparam \d_writedata[16] .is_wysiwyg = "true";
defparam \d_writedata[16] .power_up = "low";

dffeas \d_writedata[17] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[17]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_17),
	.prn(vcc));
defparam \d_writedata[17] .is_wysiwyg = "true";
defparam \d_writedata[17] .power_up = "low";

dffeas \d_writedata[18] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[18]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_18),
	.prn(vcc));
defparam \d_writedata[18] .is_wysiwyg = "true";
defparam \d_writedata[18] .power_up = "low";

dffeas \d_writedata[19] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[19]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_19),
	.prn(vcc));
defparam \d_writedata[19] .is_wysiwyg = "true";
defparam \d_writedata[19] .power_up = "low";

dffeas \d_writedata[20] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[20]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_20),
	.prn(vcc));
defparam \d_writedata[20] .is_wysiwyg = "true";
defparam \d_writedata[20] .power_up = "low";

dffeas \d_writedata[21] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[21]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_21),
	.prn(vcc));
defparam \d_writedata[21] .is_wysiwyg = "true";
defparam \d_writedata[21] .power_up = "low";

dffeas \d_writedata[22] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[22]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_22),
	.prn(vcc));
defparam \d_writedata[22] .is_wysiwyg = "true";
defparam \d_writedata[22] .power_up = "low";

dffeas \d_writedata[23] (
	.clk(wire_pll7_clk_0),
	.d(\E_st_data[23]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_23),
	.prn(vcc));
defparam \d_writedata[23] .is_wysiwyg = "true";
defparam \d_writedata[23] .power_up = "low";

cycloneive_lcell_comb \F_iw[0]~5 (
	.dataa(mem_54_0),
	.datab(data_reg_0),
	.datac(out_payload_0),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(F_iw_0),
	.cout());
defparam \F_iw[0]~5 .lut_mask = 16'hFEFF;
defparam \F_iw[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[2]~10 (
	.dataa(mem_54_0),
	.datab(data_reg_2),
	.datac(out_payload_2),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(F_iw_2),
	.cout());
defparam \F_iw[2]~10 .lut_mask = 16'hFEFF;
defparam \F_iw[2]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[12]~23 (
	.dataa(mem_54_0),
	.datab(data_reg_12),
	.datac(out_payload_12),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(F_iw_12),
	.cout());
defparam \F_iw[12]~23 .lut_mask = 16'hFEFF;
defparam \F_iw[12]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~28 (
	.dataa(mem_54_0),
	.datab(data_reg_14),
	.datac(out_payload_14),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(F_iw_14),
	.cout());
defparam \F_iw[14]~28 .lut_mask = 16'hFEFF;
defparam \F_iw[14]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[10]~33 (
	.dataa(mem_54_0),
	.datab(data_reg_10),
	.datac(out_payload_10),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(F_iw_10),
	.cout());
defparam \F_iw[10]~33 .lut_mask = 16'hFEFF;
defparam \F_iw[10]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[9]~36 (
	.dataa(mem_54_0),
	.datab(data_reg_9),
	.datac(out_payload_9),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(F_iw_9),
	.cout());
defparam \F_iw[9]~36 .lut_mask = 16'hFEFF;
defparam \F_iw[9]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[8]~39 (
	.dataa(mem_54_0),
	.datab(data_reg_8),
	.datac(out_payload_8),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(F_iw_8),
	.cout());
defparam \F_iw[8]~39 .lut_mask = 16'hFEFF;
defparam \F_iw[8]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[7]~42 (
	.dataa(mem_54_0),
	.datab(data_reg_7),
	.datac(out_payload_7),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(F_iw_7),
	.cout());
defparam \F_iw[7]~42 .lut_mask = 16'hFEFF;
defparam \F_iw[7]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~45 (
	.dataa(mem_54_0),
	.datab(data_reg_6),
	.datac(out_payload_6),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(F_iw_6),
	.cout());
defparam \F_iw[6]~45 .lut_mask = 16'hFEFF;
defparam \F_iw[6]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_valid~0 (
	.dataa(src1_valid1),
	.datab(out_valid),
	.datac(src1_valid),
	.datad(i_read1),
	.cin(gnd),
	.combout(\F_valid~0_combout ),
	.cout());
defparam \F_valid~0 .lut_mask = 16'hFEFF;
defparam \F_valid~0 .sum_lutc_input = "datac";

dffeas D_valid(
	.clk(wire_pll7_clk_0),
	.d(\F_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_valid~q ),
	.prn(vcc));
defparam D_valid.is_wysiwyg = "true";
defparam D_valid.power_up = "low";

dffeas R_valid(
	.clk(wire_pll7_clk_0),
	.d(\D_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_valid~q ),
	.prn(vcc));
defparam R_valid.is_wysiwyg = "true";
defparam R_valid.power_up = "low";

cycloneive_lcell_comb \F_iw[11]~16 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_11),
	.datad(out_data_buffer_11),
	.cin(gnd),
	.combout(\F_iw[11]~16_combout ),
	.cout());
defparam \F_iw[11]~16 .lut_mask = 16'hFFFE;
defparam \F_iw[11]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[8]~38 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_8),
	.datad(out_data_buffer_8),
	.cin(gnd),
	.combout(\F_iw[8]~38_combout ),
	.cout());
defparam \F_iw[8]~38 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[8]~40 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[8]~38_combout ),
	.datac(src1_valid1),
	.datad(F_iw_8),
	.cin(gnd),
	.combout(\F_iw[8]~40_combout ),
	.cout());
defparam \F_iw[8]~40 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~40 .sum_lutc_input = "datac";

dffeas \D_iw[8] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[8]~40_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

cycloneive_lcell_comb \F_iw[4]~14 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_4),
	.datad(out_data_buffer_4),
	.cin(gnd),
	.combout(\F_iw[4]~14_combout ),
	.cout());
defparam \F_iw[4]~14 .lut_mask = 16'hFFFE;
defparam \F_iw[4]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[4]~15 (
	.dataa(\F_iw[4]~14_combout ),
	.datab(src1_valid1),
	.datac(src_data_4),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[4]~15_combout ),
	.cout());
defparam \F_iw[4]~15 .lut_mask = 16'hFEFF;
defparam \F_iw[4]~15 .sum_lutc_input = "datac";

dffeas \D_iw[4] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[4]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

cycloneive_lcell_comb \F_iw[5]~25 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_5),
	.datad(out_data_buffer_5),
	.cin(gnd),
	.combout(\F_iw[5]~25_combout ),
	.cout());
defparam \F_iw[5]~25 .lut_mask = 16'hFFFE;
defparam \F_iw[5]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[5]~26 (
	.dataa(\F_iw[5]~25_combout ),
	.datab(src1_valid1),
	.datac(src_data_5),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[5]~26_combout ),
	.cout());
defparam \F_iw[5]~26 .lut_mask = 16'hFEFF;
defparam \F_iw[5]~26 .sum_lutc_input = "datac";

dffeas \D_iw[5] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[5]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

cycloneive_lcell_comb \F_iw[0]~4 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_0),
	.datad(out_data_buffer_0),
	.cin(gnd),
	.combout(\F_iw[0]~4_combout ),
	.cout());
defparam \F_iw[0]~4 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[0]~6 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[0]~4_combout ),
	.datac(src1_valid1),
	.datad(F_iw_0),
	.cin(gnd),
	.combout(\F_iw[0]~6_combout ),
	.cout());
defparam \F_iw[0]~6 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~6 .sum_lutc_input = "datac";

dffeas \D_iw[0] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[0]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

cycloneive_lcell_comb \F_iw[1]~7 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_1),
	.datad(out_data_buffer_1),
	.cin(gnd),
	.combout(\F_iw[1]~7_combout ),
	.cout());
defparam \F_iw[1]~7 .lut_mask = 16'hFFFE;
defparam \F_iw[1]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[1]~8 (
	.dataa(\F_iw[1]~7_combout ),
	.datab(src1_valid1),
	.datac(src_data_1),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[1]~8_combout ),
	.cout());
defparam \F_iw[1]~8 .lut_mask = 16'hFEFF;
defparam \F_iw[1]~8 .sum_lutc_input = "datac";

dffeas \D_iw[1] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[1]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

cycloneive_lcell_comb \F_iw[3]~12 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_3),
	.datad(out_data_buffer_3),
	.cin(gnd),
	.combout(\F_iw[3]~12_combout ),
	.cout());
defparam \F_iw[3]~12 .lut_mask = 16'hFFFE;
defparam \F_iw[3]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[3]~13 (
	.dataa(\F_iw[3]~12_combout ),
	.datab(src1_valid1),
	.datac(src_data_3),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[3]~13_combout ),
	.cout());
defparam \F_iw[3]~13 .lut_mask = 16'hFEFF;
defparam \F_iw[3]~13 .sum_lutc_input = "datac";

dffeas \D_iw[3] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[3]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

cycloneive_lcell_comb \F_iw[2]~9 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_2),
	.datad(out_data_buffer_2),
	.cin(gnd),
	.combout(\F_iw[2]~9_combout ),
	.cout());
defparam \F_iw[2]~9 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[2]~11 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[2]~9_combout ),
	.datac(src1_valid1),
	.datad(F_iw_2),
	.cin(gnd),
	.combout(\F_iw[2]~11_combout ),
	.cout());
defparam \F_iw[2]~11 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~11 .sum_lutc_input = "datac";

dffeas \D_iw[2] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[2]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

cycloneive_lcell_comb \Equal0~7 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
defparam \Equal0~7 .lut_mask = 16'hEFEF;
defparam \Equal0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~8 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\D_iw[0]~q ),
	.datad(\Equal0~7_combout ),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
defparam \Equal0~8 .lut_mask = 16'hFFEF;
defparam \Equal0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[15]~30 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_15),
	.datad(out_data_buffer_15),
	.cin(gnd),
	.combout(\F_iw[15]~30_combout ),
	.cout());
defparam \F_iw[15]~30 .lut_mask = 16'hFFFE;
defparam \F_iw[15]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[15]~31 (
	.dataa(\F_iw[15]~30_combout ),
	.datab(src1_valid1),
	.datac(src_data_15),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[15]~31_combout ),
	.cout());
defparam \F_iw[15]~31 .lut_mask = 16'hFEFF;
defparam \F_iw[15]~31 .sum_lutc_input = "datac";

dffeas \D_iw[15] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[15]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

dffeas E_new_inst(
	.clk(wire_pll7_clk_0),
	.d(\R_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_new_inst~q ),
	.prn(vcc));
defparam E_new_inst.is_wysiwyg = "true";
defparam E_new_inst.power_up = "low";

cycloneive_lcell_comb \D_ctrl_st~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_st~0_combout ),
	.cout());
defparam \D_ctrl_st~0 .lut_mask = 16'hBFFF;
defparam \D_ctrl_st~0 .sum_lutc_input = "datac";

dffeas R_ctrl_st(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\D_iw[2]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_st~q ),
	.prn(vcc));
defparam R_ctrl_st.is_wysiwyg = "true";
defparam R_ctrl_st.power_up = "low";

cycloneive_lcell_comb \W_valid~3 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_st~q ),
	.datac(\E_valid_from_R~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_valid~3_combout ),
	.cout());
defparam \W_valid~3 .lut_mask = 16'hF7F7;
defparam \W_valid~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_valid~2 (
	.dataa(\E_stall~4_combout ),
	.datab(d_write1),
	.datac(av_waitrequest),
	.datad(\W_valid~3_combout ),
	.cin(gnd),
	.combout(\W_valid~2_combout ),
	.cout());
defparam \W_valid~2 .lut_mask = 16'hFF7F;
defparam \W_valid~2 .sum_lutc_input = "datac";

dffeas W_valid(
	.clk(wire_pll7_clk_0),
	.d(\W_valid~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_valid~q ),
	.prn(vcc));
defparam W_valid.is_wysiwyg = "true";
defparam W_valid.power_up = "low";

cycloneive_lcell_comb \hbreak_pending_nxt~0 (
	.dataa(\hbreak_pending~q ),
	.datab(\hbreak_req~0_combout ),
	.datac(gnd),
	.datad(hbreak_enabled1),
	.cin(gnd),
	.combout(\hbreak_pending_nxt~0_combout ),
	.cout());
defparam \hbreak_pending_nxt~0 .lut_mask = 16'hEEFF;
defparam \hbreak_pending_nxt~0 .sum_lutc_input = "datac";

dffeas hbreak_pending(
	.clk(wire_pll7_clk_0),
	.d(\hbreak_pending_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\hbreak_pending~q ),
	.prn(vcc));
defparam hbreak_pending.is_wysiwyg = "true";
defparam hbreak_pending.power_up = "low";

cycloneive_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datab(hbreak_enabled1),
	.datac(\wait_for_one_post_bret_inst~q ),
	.datad(\F_valid~0_combout ),
	.cin(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.cout());
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 16'hFEFF;
defparam \wait_for_one_post_bret_inst~0 .sum_lutc_input = "datac";

dffeas wait_for_one_post_bret_inst(
	.clk(wire_pll7_clk_0),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cycloneive_lcell_comb \hbreak_req~0 (
	.dataa(\W_valid~q ),
	.datab(\hbreak_pending~q ),
	.datac(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_oci_debug|jtag_break~q ),
	.datad(\wait_for_one_post_bret_inst~q ),
	.cin(gnd),
	.combout(\hbreak_req~0_combout ),
	.cout());
defparam \hbreak_req~0 .lut_mask = 16'hFEFF;
defparam \hbreak_req~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~27 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_14),
	.datad(out_data_buffer_14),
	.cin(gnd),
	.combout(\F_iw[14]~27_combout ),
	.cout());
defparam \F_iw[14]~27 .lut_mask = 16'hFFFE;
defparam \F_iw[14]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~29 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[14]~27_combout ),
	.datac(src1_valid1),
	.datad(F_iw_14),
	.cin(gnd),
	.combout(\F_iw[14]~29_combout ),
	.cout());
defparam \F_iw[14]~29 .lut_mask = 16'hFFFE;
defparam \F_iw[14]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~78 (
	.dataa(\D_iw[1]~1_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\F_iw[14]~29_combout ),
	.cin(gnd),
	.combout(\F_iw[14]~78_combout ),
	.cout());
defparam \F_iw[14]~78 .lut_mask = 16'hFFDF;
defparam \F_iw[14]~78 .sum_lutc_input = "datac";

dffeas \D_iw[14] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[14]~78_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

cycloneive_lcell_comb \D_op_opx_rsv63~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_op_opx_rsv63~0_combout ),
	.cout());
defparam \D_op_opx_rsv63~0 .lut_mask = 16'hEEEE;
defparam \D_op_opx_rsv63~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[13]~18 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_13),
	.datad(out_data_buffer_13),
	.cin(gnd),
	.combout(\F_iw[13]~18_combout ),
	.cout());
defparam \F_iw[13]~18 .lut_mask = 16'hFFFE;
defparam \F_iw[13]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[13]~19 (
	.dataa(\F_iw[13]~18_combout ),
	.datab(src1_valid1),
	.datac(src_data_13),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[13]~19_combout ),
	.cout());
defparam \F_iw[13]~19 .lut_mask = 16'hFEFF;
defparam \F_iw[13]~19 .sum_lutc_input = "datac";

dffeas \D_iw[13] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[13]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

cycloneive_lcell_comb \F_iw[16]~20 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_16),
	.datad(out_data_buffer_16),
	.cin(gnd),
	.combout(\F_iw[16]~20_combout ),
	.cout());
defparam \F_iw[16]~20 .lut_mask = 16'hFFFE;
defparam \F_iw[16]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[16]~21 (
	.dataa(\F_iw[16]~20_combout ),
	.datab(out_payload_0),
	.datac(src_payload),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[16]~21_combout ),
	.cout());
defparam \F_iw[16]~21 .lut_mask = 16'hFEFF;
defparam \F_iw[16]~21 .sum_lutc_input = "datac";

dffeas \D_iw[16] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[16]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

cycloneive_lcell_comb \F_iw[12]~22 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_12),
	.datad(out_data_buffer_12),
	.cin(gnd),
	.combout(\F_iw[12]~22_combout ),
	.cout());
defparam \F_iw[12]~22 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[12]~24 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[12]~22_combout ),
	.datac(src1_valid1),
	.datad(F_iw_12),
	.cin(gnd),
	.combout(\F_iw[12]~24_combout ),
	.cout());
defparam \F_iw[12]~24 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~24 .sum_lutc_input = "datac";

dffeas \D_iw[12] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[12]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

cycloneive_lcell_comb \Equal62~4 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~4_combout ),
	.cout());
defparam \Equal62~4 .lut_mask = 16'hFF7F;
defparam \Equal62~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~5 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~5_combout ),
	.cout());
defparam \Equal62~5 .lut_mask = 16'hFFF7;
defparam \Equal62~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~6 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~6_combout ),
	.cout());
defparam \Equal62~6 .lut_mask = 16'hFFFB;
defparam \Equal62~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~4_combout ),
	.datac(\Equal62~5_combout ),
	.datad(\Equal62~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_shift_rot~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~7 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~7_combout ),
	.cout());
defparam \Equal62~7 .lut_mask = 16'hFFBF;
defparam \Equal62~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(\Equal62~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot~1 .lut_mask = 16'hEEFF;
defparam \D_ctrl_shift_rot~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_logical~0 (
	.dataa(\D_iw[12]~q ),
	.datab(gnd),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~0_combout ),
	.cout());
defparam \D_ctrl_shift_logical~0 .lut_mask = 16'hAFFF;
defparam \D_ctrl_shift_logical~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~2 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\Equal62~4_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~2_combout ),
	.cout());
defparam \D_ctrl_shift_rot~2 .lut_mask = 16'hACFF;
defparam \D_ctrl_shift_rot~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~3 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_ctrl_shift_rot~0_combout ),
	.datac(\D_ctrl_shift_rot~1_combout ),
	.datad(\D_ctrl_shift_rot~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~3_combout ),
	.cout());
defparam \D_ctrl_shift_rot~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_shift_rot~3 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_shift_rot~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_shift_rot.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[0]~5 (
	.dataa(\E_shift_rot_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\E_shift_rot_cnt[0]~5_combout ),
	.cout(\E_shift_rot_cnt[0]~6 ));
defparam \E_shift_rot_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \E_shift_rot_cnt[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_hi_imm16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~0_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~0 .lut_mask = 16'hFFF7;
defparam \D_ctrl_hi_imm16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_hi_imm16~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\D_ctrl_hi_imm16~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~1_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~1 .lut_mask = 16'hFEFE;
defparam \D_ctrl_hi_imm16~1 .sum_lutc_input = "datac";

dffeas R_ctrl_hi_imm16(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_hi_imm16~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam R_ctrl_hi_imm16.is_wysiwyg = "true";
defparam R_ctrl_hi_imm16.power_up = "low";

cycloneive_lcell_comb \Equal0~14 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~14_combout ),
	.cout());
defparam \Equal0~14 .lut_mask = 16'hDFFF;
defparam \Equal0~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~14 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[0]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~14_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~14 .lut_mask = 16'hF6FF;
defparam \D_ctrl_alu_force_xor~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~15 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~15_combout ),
	.cout());
defparam \Equal0~15 .lut_mask = 16'hFFFE;
defparam \Equal0~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~16 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~16_combout ),
	.cout());
defparam \Equal0~16 .lut_mask = 16'hFFFD;
defparam \Equal0~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~0 (
	.dataa(\D_iw[5]~q ),
	.datab(\D_ctrl_alu_force_xor~14_combout ),
	.datac(\Equal0~15_combout ),
	.datad(\Equal0~16_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~0_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~0 .lut_mask = 16'h7FFF;
defparam \D_ctrl_force_src2_zero~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~14 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~14_combout ),
	.cout());
defparam \Equal62~14 .lut_mask = 16'hFEFF;
defparam \Equal62~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~13 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~13_combout ),
	.cout());
defparam \Equal62~13 .lut_mask = 16'hFDFF;
defparam \Equal62~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~1 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~14_combout ),
	.datac(\Equal62~13_combout ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~1_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~8 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~8_combout ),
	.cout());
defparam \Equal62~8 .lut_mask = 16'hEFFF;
defparam \Equal62~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~2 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_ctrl_force_src2_zero~1_combout ),
	.datac(\Equal62~8_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~2_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~2 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~13 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~13_combout ),
	.cout());
defparam \Equal0~13 .lut_mask = 16'hBFFF;
defparam \Equal0~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFBFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~3 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~13_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~3_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~3 .lut_mask = 16'hFFDE;
defparam \D_ctrl_force_src2_zero~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~4 (
	.dataa(\D_ctrl_force_src2_zero~0_combout ),
	.datab(\D_ctrl_force_src2_zero~2_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_force_src2_zero~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~4_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~4 .lut_mask = 16'hFFFD;
defparam \D_ctrl_force_src2_zero~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~9 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~9_combout ),
	.cout());
defparam \Equal62~9 .lut_mask = 16'hBFFF;
defparam \Equal62~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~1 (
	.dataa(\D_iw[15]~q ),
	.datab(gnd),
	.datac(\Equal0~8_combout ),
	.datad(\Equal62~9_combout ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~1_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~1 .lut_mask = 16'hAFFF;
defparam \D_ctrl_uncond_cti_non_br~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~10 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~10_combout ),
	.cout());
defparam \Equal62~10 .lut_mask = 16'hFFEF;
defparam \Equal62~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hEEEE;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_cmpge~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_cmpge~0_combout ),
	.cout());
defparam \D_op_cmpge~0 .lut_mask = 16'hFEFF;
defparam \D_op_cmpge~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~13 (
	.dataa(gnd),
	.datab(\Equal62~4_combout ),
	.datac(\Equal62~10_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~13_combout ),
	.cout());
defparam \D_ctrl_exception~13 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~11 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~11_combout ),
	.cout());
defparam \Equal62~11 .lut_mask = 16'hDFFF;
defparam \Equal62~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_opx_rsv17~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv17~0_combout ),
	.cout());
defparam \D_op_opx_rsv17~0 .lut_mask = 16'hFEFF;
defparam \D_op_opx_rsv17~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~14 (
	.dataa(gnd),
	.datab(\Equal62~9_combout ),
	.datac(\Equal62~11_combout ),
	.datad(\D_op_opx_rsv17~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~14_combout ),
	.cout());
defparam \D_ctrl_exception~14 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~2 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~2_combout ),
	.cout());
defparam \Equal62~2 .lut_mask = 16'hFBFF;
defparam \Equal62~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_opx_rsv00~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~2_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv00~0_combout ),
	.cout());
defparam \D_op_opx_rsv00~0 .lut_mask = 16'hFEFF;
defparam \D_op_opx_rsv00~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~15 (
	.dataa(\D_iw[14]~q ),
	.datab(\Equal62~2_combout ),
	.datac(\Equal62~0_combout ),
	.datad(\D_op_opx_rsv00~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~15_combout ),
	.cout());
defparam \D_ctrl_exception~15 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~16 (
	.dataa(\D_iw[14]~q ),
	.datab(\Equal62~5_combout ),
	.datac(\Equal62~6_combout ),
	.datad(\D_op_opx_rsv00~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~16_combout ),
	.cout());
defparam \D_ctrl_exception~16 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~17 (
	.dataa(\D_ctrl_exception~13_combout ),
	.datab(\D_ctrl_exception~14_combout ),
	.datac(\D_ctrl_exception~15_combout ),
	.datad(\D_ctrl_exception~16_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~17_combout ),
	.cout());
defparam \D_ctrl_exception~17 .lut_mask = 16'hFFFE;
defparam \D_ctrl_exception~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~18 (
	.dataa(\Equal62~6_combout ),
	.datab(\D_op_opx_rsv17~0_combout ),
	.datac(\Equal62~5_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~18_combout ),
	.cout());
defparam \D_ctrl_exception~18 .lut_mask = 16'h7FFF;
defparam \D_ctrl_exception~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~12 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~12_combout ),
	.cout());
defparam \Equal0~12 .lut_mask = 16'hFDFF;
defparam \Equal0~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~19 (
	.dataa(\D_op_opx_rsv17~0_combout ),
	.datab(\Equal0~12_combout ),
	.datac(\Equal62~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_exception~19_combout ),
	.cout());
defparam \D_ctrl_exception~19 .lut_mask = 16'h7F7F;
defparam \D_ctrl_exception~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~12 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~12_combout ),
	.cout());
defparam \Equal62~12 .lut_mask = 16'hFFFE;
defparam \Equal62~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~3 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~3_combout ),
	.cout());
defparam \Equal62~3 .lut_mask = 16'hFFFD;
defparam \Equal62~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~1 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~1_combout ),
	.cout());
defparam \Equal62~1 .lut_mask = 16'hF7FF;
defparam \Equal62~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~20 (
	.dataa(\Equal62~3_combout ),
	.datab(\Equal62~13_combout ),
	.datac(\Equal62~1_combout ),
	.datad(\Equal62~9_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~20_combout ),
	.cout());
defparam \D_ctrl_exception~20 .lut_mask = 16'h7FFF;
defparam \D_ctrl_exception~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~23 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~12_combout ),
	.datad(\D_ctrl_exception~20_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~23_combout ),
	.cout());
defparam \D_ctrl_exception~23 .lut_mask = 16'hFF7F;
defparam \D_ctrl_exception~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~21 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_ctrl_exception~18_combout ),
	.datac(\D_ctrl_exception~19_combout ),
	.datad(\D_ctrl_exception~23_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~21_combout ),
	.cout());
defparam \D_ctrl_exception~21 .lut_mask = 16'hFFFD;
defparam \D_ctrl_exception~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'h7FFF;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_jmp_direct~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~0_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~0 .lut_mask = 16'h0FFF;
defparam \D_ctrl_jmp_direct~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~11_combout ),
	.datac(\Equal62~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.cout());
defparam \D_ctrl_retaddr~0 .lut_mask = 16'hFEFE;
defparam \D_ctrl_retaddr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(\Equal62~14_combout ),
	.datab(\Equal62~13_combout ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.cout());
defparam \D_ctrl_retaddr~1 .lut_mask = 16'hEEFF;
defparam \D_ctrl_retaddr~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~2 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_retaddr~0_combout ),
	.datad(\D_ctrl_retaddr~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~2_combout ),
	.cout());
defparam \D_ctrl_retaddr~2 .lut_mask = 16'hFFFE;
defparam \D_ctrl_retaddr~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~5 (
	.dataa(\Equal0~4_combout ),
	.datab(\Equal0~13_combout ),
	.datac(\D_ctrl_jmp_direct~0_combout ),
	.datad(\D_ctrl_retaddr~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~5_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~5 .lut_mask = 16'h7FFF;
defparam \D_ctrl_force_src2_zero~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~18 (
	.dataa(\Equal0~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\Equal0~18_combout ),
	.cout());
defparam \Equal0~18 .lut_mask = 16'hAAFF;
defparam \Equal0~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~6 (
	.dataa(\D_ctrl_exception~17_combout ),
	.datab(\D_ctrl_exception~21_combout ),
	.datac(\D_ctrl_force_src2_zero~5_combout ),
	.datad(\Equal0~18_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~6_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~6 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~7 (
	.dataa(\Equal0~14_combout ),
	.datab(\D_ctrl_force_src2_zero~4_combout ),
	.datac(\D_ctrl_uncond_cti_non_br~1_combout ),
	.datad(\D_ctrl_force_src2_zero~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~7_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~7 .lut_mask = 16'hEFFF;
defparam \D_ctrl_force_src2_zero~7 .sum_lutc_input = "datac";

dffeas R_ctrl_force_src2_zero(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_force_src2_zero~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_force_src2_zero~q ),
	.prn(vcc));
defparam R_ctrl_force_src2_zero.is_wysiwyg = "true";
defparam R_ctrl_force_src2_zero.power_up = "low";

cycloneive_lcell_comb \R_src2_lo[4]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\R_ctrl_hi_imm16~q ),
	.datad(\R_ctrl_force_src2_zero~q ),
	.cin(gnd),
	.combout(\R_src2_lo[4]~2_combout ),
	.cout());
defparam \R_src2_lo[4]~2 .lut_mask = 16'h0FFF;
defparam \R_src2_lo[4]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~44 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_6),
	.datad(out_data_buffer_6),
	.cin(gnd),
	.combout(\F_iw[6]~44_combout ),
	.cout());
defparam \F_iw[6]~44 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~46 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[6]~44_combout ),
	.datac(src1_valid1),
	.datad(F_iw_6),
	.cin(gnd),
	.combout(\F_iw[6]~46_combout ),
	.cout());
defparam \F_iw[6]~46 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~46 .sum_lutc_input = "datac";

dffeas \D_iw[6] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[6]~46_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

cycloneive_lcell_comb \D_ctrl_src_imm5_shift_rot~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~0 .lut_mask = 16'hBBF3;
defparam \D_ctrl_src_imm5_shift_rot~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_src_imm5_shift_rot~1 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~1 .lut_mask = 16'hEFFF;
defparam \D_ctrl_src_imm5_shift_rot~1 .sum_lutc_input = "datac";

dffeas R_ctrl_src_imm5_shift_rot(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_src_imm5_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_src_imm5_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_src_imm5_shift_rot.power_up = "low";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~7 (
	.dataa(\D_iw[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~7_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~7 .lut_mask = 16'hAAFF;
defparam \D_ctrl_implicit_dst_eretaddr~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~0 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~5_combout ),
	.datac(\Equal62~4_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~0_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_unsigned_lo_imm16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~1 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_ctrl_unsigned_lo_imm16~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~1_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~1 .lut_mask = 16'hEEEE;
defparam \D_ctrl_unsigned_lo_imm16~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~17 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~17_combout ),
	.cout());
defparam \Equal0~17 .lut_mask = 16'hFFDF;
defparam \Equal0~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~0 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~0_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~0 .lut_mask = 16'h6996;
defparam \D_ctrl_b_is_dst~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~1_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~1 .lut_mask = 16'hFBFE;
defparam \D_ctrl_b_is_dst~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~2 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_ctrl_b_is_dst~0_combout ),
	.datad(\D_ctrl_b_is_dst~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~2_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~2 .lut_mask = 16'h96FF;
defparam \D_ctrl_b_is_dst~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_use_imm~0 (
	.dataa(\Equal0~17_combout ),
	.datab(\D_ctrl_b_is_dst~2_combout ),
	.datac(\Equal0~16_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\R_src2_use_imm~0_combout ),
	.cout());
defparam \R_src2_use_imm~0 .lut_mask = 16'hFEFF;
defparam \R_src2_use_imm~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_ctrl_br_nxt~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[4]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~0_combout ),
	.cout());
defparam \R_ctrl_br_nxt~0 .lut_mask = 16'hFFFE;
defparam \R_ctrl_br_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_ctrl_br_nxt~1 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_br_nxt~0_combout ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~1_combout ),
	.cout());
defparam \R_ctrl_br_nxt~1 .lut_mask = 16'hEEFF;
defparam \R_ctrl_br_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_use_imm~1 (
	.dataa(\D_ctrl_unsigned_lo_imm16~1_combout ),
	.datab(\R_src2_use_imm~0_combout ),
	.datac(\R_valid~q ),
	.datad(\R_ctrl_br_nxt~1_combout ),
	.cin(gnd),
	.combout(\R_src2_use_imm~1_combout ),
	.cout());
defparam \R_src2_use_imm~1 .lut_mask = 16'hFFFE;
defparam \R_src2_use_imm~1 .sum_lutc_input = "datac";

dffeas R_src2_use_imm(
	.clk(wire_pll7_clk_0),
	.d(\R_src2_use_imm~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_src2_use_imm~q ),
	.prn(vcc));
defparam R_src2_use_imm.is_wysiwyg = "true";
defparam R_src2_use_imm.power_up = "low";

cycloneive_lcell_comb \R_src2_lo~3 (
	.dataa(\R_ctrl_src_imm5_shift_rot~q ),
	.datab(\R_src2_use_imm~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\R_src2_lo~3_combout ),
	.cout());
defparam \R_src2_lo~3 .lut_mask = 16'hEEEE;
defparam \R_src2_lo~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[0]~8 (
	.dataa(\R_src2_lo[4]~2_combout ),
	.datab(\D_iw[6]~q ),
	.datac(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\R_src2_lo~3_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[0]~8_combout ),
	.cout());
defparam \R_src2_lo[0]~8 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[0]~8 .sum_lutc_input = "datac";

dffeas \E_src2[0] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

dffeas \E_shift_rot_cnt[0] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_cnt[0]~5_combout ),
	.asdata(\E_src2[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[0] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[0] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[1]~7 (
	.dataa(\E_shift_rot_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[0]~6 ),
	.combout(\E_shift_rot_cnt[1]~7_combout ),
	.cout(\E_shift_rot_cnt[1]~8 ));
defparam \E_shift_rot_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[1]~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[7]~41 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_7),
	.datad(out_data_buffer_7),
	.cin(gnd),
	.combout(\F_iw[7]~41_combout ),
	.cout());
defparam \F_iw[7]~41 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[7]~43 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[7]~41_combout ),
	.datac(src1_valid1),
	.datad(F_iw_7),
	.cin(gnd),
	.combout(\F_iw[7]~43_combout ),
	.cout());
defparam \F_iw[7]~43 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~43 .sum_lutc_input = "datac";

dffeas \D_iw[7] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[7]~43_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[1]~7 (
	.dataa(\R_src2_lo[4]~2_combout ),
	.datab(\D_iw[7]~q ),
	.datac(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\R_src2_lo~3_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[1]~7_combout ),
	.cout());
defparam \R_src2_lo[1]~7 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[1]~7 .sum_lutc_input = "datac";

dffeas \E_src2[1] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[1]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

dffeas \E_shift_rot_cnt[1] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_cnt[1]~7_combout ),
	.asdata(\E_src2[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[1] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[1] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[2]~9 (
	.dataa(\E_shift_rot_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[1]~8 ),
	.combout(\E_shift_rot_cnt[2]~9_combout ),
	.cout(\E_shift_rot_cnt[2]~10 ));
defparam \E_shift_rot_cnt[2]~9 .lut_mask = 16'h5AAF;
defparam \E_shift_rot_cnt[2]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \R_src2_lo[2]~6 (
	.dataa(\R_src2_lo[4]~2_combout ),
	.datab(\D_iw[8]~q ),
	.datac(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datad(\R_src2_lo~3_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[2]~6_combout ),
	.cout());
defparam \R_src2_lo[2]~6 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[2]~6 .sum_lutc_input = "datac";

dffeas \E_src2[2] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[2]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

dffeas \E_shift_rot_cnt[2] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_cnt[2]~9_combout ),
	.asdata(\E_src2[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[2] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[2] .power_up = "low";

cycloneive_lcell_comb \E_stall~0 (
	.dataa(\E_new_inst~q ),
	.datab(\E_shift_rot_cnt[0]~q ),
	.datac(\E_shift_rot_cnt[1]~q ),
	.datad(\E_shift_rot_cnt[2]~q ),
	.cin(gnd),
	.combout(\E_stall~0_combout ),
	.cout());
defparam \E_stall~0 .lut_mask = 16'hFFFE;
defparam \E_stall~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_shift_rot_cnt[3]~11 (
	.dataa(\E_shift_rot_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[2]~10 ),
	.combout(\E_shift_rot_cnt[3]~11_combout ),
	.cout(\E_shift_rot_cnt[3]~12 ));
defparam \E_shift_rot_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[3]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[9]~35 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_9),
	.datad(out_data_buffer_9),
	.cin(gnd),
	.combout(\F_iw[9]~35_combout ),
	.cout());
defparam \F_iw[9]~35 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[9]~37 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[9]~35_combout ),
	.datac(src1_valid1),
	.datad(F_iw_9),
	.cin(gnd),
	.combout(\F_iw[9]~37_combout ),
	.cout());
defparam \F_iw[9]~37 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~37 .sum_lutc_input = "datac";

dffeas \D_iw[9] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[9]~37_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[3]~5 (
	.dataa(\R_src2_lo[4]~2_combout ),
	.datab(\D_iw[9]~q ),
	.datac(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datad(\R_src2_lo~3_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[3]~5_combout ),
	.cout());
defparam \R_src2_lo[3]~5 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[3]~5 .sum_lutc_input = "datac";

dffeas \E_src2[3] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

dffeas \E_shift_rot_cnt[3] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_cnt[3]~11_combout ),
	.asdata(\E_src2[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[3] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[3] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[4]~13 (
	.dataa(\E_shift_rot_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\E_shift_rot_cnt[3]~12 ),
	.combout(\E_shift_rot_cnt[4]~13_combout ),
	.cout());
defparam \E_shift_rot_cnt[4]~13 .lut_mask = 16'h5A5A;
defparam \E_shift_rot_cnt[4]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[10]~32 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_10),
	.datad(out_data_buffer_10),
	.cin(gnd),
	.combout(\F_iw[10]~32_combout ),
	.cout());
defparam \F_iw[10]~32 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[10]~34 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[10]~32_combout ),
	.datac(src1_valid1),
	.datad(F_iw_10),
	.cin(gnd),
	.combout(\F_iw[10]~34_combout ),
	.cout());
defparam \F_iw[10]~34 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~34 .sum_lutc_input = "datac";

dffeas \D_iw[10] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[10]~34_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[4]~4 (
	.dataa(\R_src2_lo[4]~2_combout ),
	.datab(\D_iw[10]~q ),
	.datac(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datad(\R_src2_lo~3_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[4]~4_combout ),
	.cout());
defparam \R_src2_lo[4]~4 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[4]~4 .sum_lutc_input = "datac";

dffeas \E_src2[4] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

dffeas \E_shift_rot_cnt[4] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_cnt[4]~13_combout ),
	.asdata(\E_src2[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[4] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[4] .power_up = "low";

cycloneive_lcell_comb \E_stall~1 (
	.dataa(\E_shift_rot_cnt[3]~q ),
	.datab(\E_shift_rot_cnt[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_stall~1_combout ),
	.cout());
defparam \E_stall~1 .lut_mask = 16'hEEEE;
defparam \E_stall~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~2 (
	.dataa(\R_ctrl_shift_rot~q ),
	.datab(\E_valid_from_R~q ),
	.datac(\E_stall~0_combout ),
	.datad(\E_stall~1_combout ),
	.cin(gnd),
	.combout(\E_stall~2_combout ),
	.cout());
defparam \E_stall~2 .lut_mask = 16'hFFFE;
defparam \E_stall~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld_signed~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~0_combout ),
	.cout());
defparam \D_ctrl_ld_signed~0 .lut_mask = 16'hEFFF;
defparam \D_ctrl_ld_signed~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld~2 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld~2_combout ),
	.cout());
defparam \D_ctrl_ld~2 .lut_mask = 16'hBFBF;
defparam \D_ctrl_ld~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld~3 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(\D_iw[0]~q ),
	.datad(\D_ctrl_ld~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_ld~3_combout ),
	.cout());
defparam \D_ctrl_ld~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_ld~3 .sum_lutc_input = "datac";

dffeas R_ctrl_ld(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_ld~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld~q ),
	.prn(vcc));
defparam R_ctrl_ld.is_wysiwyg = "true";
defparam R_ctrl_ld.power_up = "low";

cycloneive_lcell_comb \av_ld_waiting_for_data_nxt~0 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_waiting_for_data_nxt~0_combout ),
	.cout());
defparam \av_ld_waiting_for_data_nxt~0 .lut_mask = 16'hEEEE;
defparam \av_ld_waiting_for_data_nxt~0 .sum_lutc_input = "datac";

dffeas av_ld_waiting_for_data(
	.clk(wire_pll7_clk_0),
	.d(\av_ld_waiting_for_data_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_waiting_for_data~q ),
	.prn(vcc));
defparam av_ld_waiting_for_data.is_wysiwyg = "true";
defparam av_ld_waiting_for_data.power_up = "low";

cycloneive_lcell_comb \av_ld_waiting_for_data_nxt~1 (
	.dataa(WideOr1),
	.datab(\av_ld_waiting_for_data_nxt~0_combout ),
	.datac(\av_ld_waiting_for_data~q ),
	.datad(d_read1),
	.cin(gnd),
	.combout(\av_ld_waiting_for_data_nxt~1_combout ),
	.cout());
defparam \av_ld_waiting_for_data_nxt~1 .lut_mask = 16'hACFF;
defparam \av_ld_waiting_for_data_nxt~1 .sum_lutc_input = "datac";

dffeas av_ld_aligning_data(
	.clk(wire_pll7_clk_0),
	.d(\av_ld_aligning_data_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_aligning_data~q ),
	.prn(vcc));
defparam av_ld_aligning_data.is_wysiwyg = "true";
defparam av_ld_aligning_data.power_up = "low";

cycloneive_lcell_comb \D_ctrl_mem16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~0_combout ),
	.cout());
defparam \D_ctrl_mem16~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_mem16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem16~1 (
	.dataa(\D_ctrl_mem16~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~1_combout ),
	.cout());
defparam \D_ctrl_mem16~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem16~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_align_cycle_nxt[0]~0 (
	.dataa(\av_ld_align_cycle[0]~q ),
	.datab(d_read1),
	.datac(gnd),
	.datad(WideOr1),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[0]~0_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[0]~0 .lut_mask = 16'hFF77;
defparam \av_ld_align_cycle_nxt[0]~0 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[0] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_align_cycle_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[0]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[0] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[0] .power_up = "low";

cycloneive_lcell_comb \av_ld_align_cycle_nxt[1]~1 (
	.dataa(WideOr1),
	.datab(d_read1),
	.datac(\av_ld_align_cycle[1]~q ),
	.datad(\av_ld_align_cycle[0]~q ),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[1]~1_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[1]~1 .lut_mask = 16'hBFFB;
defparam \av_ld_align_cycle_nxt[1]~1 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[1] (
	.clk(wire_pll7_clk_0),
	.d(\av_ld_align_cycle_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[1]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[1] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[1] .power_up = "low";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~0 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\D_ctrl_mem16~1_combout ),
	.datac(\av_ld_align_cycle[0]~q ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~0_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~0 .lut_mask = 16'hBEFF;
defparam \av_ld_aligning_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem32~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem32~0_combout ),
	.cout());
defparam \D_ctrl_mem32~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem32~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\av_ld_aligning_data~q ),
	.datad(\D_ctrl_mem32~0_combout ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~1_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~1 .lut_mask = 16'h0FFF;
defparam \av_ld_aligning_data_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~2 (
	.dataa(\av_ld_aligning_data_nxt~0_combout ),
	.datab(d_read1),
	.datac(\av_ld_aligning_data_nxt~1_combout ),
	.datad(WideOr1),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~2_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~2 .lut_mask = 16'hFEFF;
defparam \av_ld_aligning_data_nxt~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~3 (
	.dataa(\E_valid_from_R~q ),
	.datab(\av_ld_waiting_for_data_nxt~1_combout ),
	.datac(\av_ld_aligning_data_nxt~2_combout ),
	.datad(\D_ctrl_mem32~0_combout ),
	.cin(gnd),
	.combout(\E_stall~3_combout ),
	.cout());
defparam \E_stall~3 .lut_mask = 16'hFEFF;
defparam \E_stall~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~4 (
	.dataa(\E_stall~2_combout ),
	.datab(\R_ctrl_ld~q ),
	.datac(\E_new_inst~q ),
	.datad(\E_stall~3_combout ),
	.cin(gnd),
	.combout(\E_stall~4_combout ),
	.cout());
defparam \E_stall~4 .lut_mask = 16'hFFFE;
defparam \E_stall~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_valid_from_R~3 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_st~q ),
	.datac(\R_valid~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_valid_from_R~3_combout ),
	.cout());
defparam \E_valid_from_R~3 .lut_mask = 16'hFEFE;
defparam \E_valid_from_R~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_valid_from_R~2 (
	.dataa(\E_stall~4_combout ),
	.datab(d_write1),
	.datac(av_waitrequest),
	.datad(\E_valid_from_R~3_combout ),
	.cin(gnd),
	.combout(\E_valid_from_R~2_combout ),
	.cout());
defparam \E_valid_from_R~2 .lut_mask = 16'hFFFE;
defparam \E_valid_from_R~2 .sum_lutc_input = "datac";

dffeas E_valid_from_R(
	.clk(wire_pll7_clk_0),
	.d(\E_valid_from_R~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_valid_from_R~q ),
	.prn(vcc));
defparam E_valid_from_R.is_wysiwyg = "true";
defparam E_valid_from_R.power_up = "low";

cycloneive_lcell_comb \D_ctrl_jmp_direct~1 (
	.dataa(\D_ctrl_jmp_direct~0_combout ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~1_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~1 .lut_mask = 16'hBFFF;
defparam \D_ctrl_jmp_direct~1 .sum_lutc_input = "datac";

dffeas R_ctrl_jmp_direct(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_jmp_direct~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_jmp_direct~q ),
	.prn(vcc));
defparam R_ctrl_jmp_direct.is_wysiwyg = "true";
defparam R_ctrl_jmp_direct.power_up = "low";

cycloneive_lcell_comb \R_src1~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_valid_from_R~q ),
	.datad(\R_ctrl_jmp_direct~q ),
	.cin(gnd),
	.combout(\R_src1~14_combout ),
	.cout());
defparam \R_src1~14 .lut_mask = 16'h0FFF;
defparam \R_src1~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[4]~22 (
	.dataa(\D_iw[8]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[4]~22_combout ),
	.cout());
defparam \E_src1[4]~22 .lut_mask = 16'hAACC;
defparam \E_src1[4]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[0]~0 (
	.dataa(F_pc_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\F_pc_plus_one[0]~0_combout ),
	.cout(\F_pc_plus_one[0]~1 ));
defparam \F_pc_plus_one[0]~0 .lut_mask = 16'h55AA;
defparam \F_pc_plus_one[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[1]~2 (
	.dataa(F_pc_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[0]~1 ),
	.combout(\F_pc_plus_one[1]~2_combout ),
	.cout(\F_pc_plus_one[1]~3 ));
defparam \F_pc_plus_one[1]~2 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[2]~4 (
	.dataa(F_pc_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[1]~3 ),
	.combout(\F_pc_plus_one[2]~4_combout ),
	.cout(\F_pc_plus_one[2]~5 ));
defparam \F_pc_plus_one[2]~4 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[2]~4 .sum_lutc_input = "cin";

dffeas R_ctrl_br(
	.clk(wire_pll7_clk_0),
	.d(\R_ctrl_br_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br~q ),
	.prn(vcc));
defparam R_ctrl_br.is_wysiwyg = "true";
defparam R_ctrl_br.power_up = "low";

cycloneive_lcell_comb \D_ctrl_retaddr~3 (
	.dataa(\Equal62~13_combout ),
	.datab(\Equal62~12_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~3_combout ),
	.cout());
defparam \D_ctrl_retaddr~3 .lut_mask = 16'hEFFF;
defparam \D_ctrl_retaddr~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~4 (
	.dataa(\D_ctrl_retaddr~3_combout ),
	.datab(\Equal62~14_combout ),
	.datac(\Equal62~10_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~4_combout ),
	.cout());
defparam \D_ctrl_retaddr~4 .lut_mask = 16'hFEFF;
defparam \D_ctrl_retaddr~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~5 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_ctrl_retaddr~4_combout ),
	.datac(\D_ctrl_force_src2_zero~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~5_combout ),
	.cout());
defparam \D_ctrl_retaddr~5 .lut_mask = 16'hF7F7;
defparam \D_ctrl_retaddr~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~10 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~10_combout ),
	.cout());
defparam \Equal0~10 .lut_mask = 16'hFF7F;
defparam \Equal0~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~6 (
	.dataa(\Equal0~14_combout ),
	.datab(\D_ctrl_force_src2_zero~0_combout ),
	.datac(\Equal0~10_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~6_combout ),
	.cout());
defparam \D_ctrl_retaddr~6 .lut_mask = 16'hFDFE;
defparam \D_ctrl_retaddr~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~7 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~13_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~7_combout ),
	.cout());
defparam \D_ctrl_retaddr~7 .lut_mask = 16'hFFBE;
defparam \D_ctrl_retaddr~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~8 (
	.dataa(\Equal0~2_combout ),
	.datab(\D_ctrl_retaddr~5_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~8_combout ),
	.cout());
defparam \D_ctrl_retaddr~8 .lut_mask = 16'hBFFB;
defparam \D_ctrl_retaddr~8 .sum_lutc_input = "datac";

dffeas R_ctrl_retaddr(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_retaddr~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_retaddr~q ),
	.prn(vcc));
defparam R_ctrl_retaddr.is_wysiwyg = "true";
defparam R_ctrl_retaddr.power_up = "low";

cycloneive_lcell_comb \R_src1~15 (
	.dataa(\R_ctrl_br~q ),
	.datab(\R_valid~q ),
	.datac(\R_ctrl_retaddr~q ),
	.datad(\E_valid_from_R~q ),
	.cin(gnd),
	.combout(\R_src1~15_combout ),
	.cout());
defparam \R_src1~15 .lut_mask = 16'hFFFE;
defparam \R_src1~15 .sum_lutc_input = "datac";

dffeas \E_src1[4] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[4]~22_combout ),
	.asdata(\F_pc_plus_one[2]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

cycloneive_lcell_comb \Equal135~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[9]~q ),
	.datad(\D_iw[10]~q ),
	.cin(gnd),
	.combout(\Equal135~0_combout ),
	.cout());
defparam \Equal135~0 .lut_mask = 16'h0FFF;
defparam \Equal135~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal135~1 (
	.dataa(\D_iw[7]~q ),
	.datab(\D_iw[6]~q ),
	.datac(\Equal135~0_combout ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\Equal135~1_combout ),
	.cout());
defparam \Equal135~1 .lut_mask = 16'hFEFF;
defparam \Equal135~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb D_op_wrctl(
	.dataa(\Equal0~8_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~3_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_wrctl~combout ),
	.cout());
defparam D_op_wrctl.lut_mask = 16'hFEFF;
defparam D_op_wrctl.sum_lutc_input = "datac";

dffeas R_ctrl_wrctl_inst(
	.clk(wire_pll7_clk_0),
	.d(\D_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam R_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam R_ctrl_wrctl_inst.power_up = "low";

cycloneive_lcell_comb \W_ienable_reg_nxt~0 (
	.dataa(\E_valid_from_R~q ),
	.datab(\Equal135~1_combout ),
	.datac(\R_ctrl_wrctl_inst~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_ienable_reg_nxt~0_combout ),
	.cout());
defparam \W_ienable_reg_nxt~0 .lut_mask = 16'hFEFE;
defparam \W_ienable_reg_nxt~0 .sum_lutc_input = "datac";

dffeas \W_ienable_reg[4] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~0_combout ),
	.q(\W_ienable_reg[4]~q ),
	.prn(vcc));
defparam \W_ienable_reg[4] .is_wysiwyg = "true";
defparam \W_ienable_reg[4] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[4]~0 (
	.dataa(\W_ienable_reg[4]~q ),
	.datab(irq),
	.datac(gnd),
	.datad(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[4]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[4]~0_combout ),
	.cout());
defparam \W_ipending_reg_nxt[4]~0 .lut_mask = 16'hEEFF;
defparam \W_ipending_reg_nxt[4]~0 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[4] (
	.clk(wire_pll7_clk_0),
	.d(\W_ipending_reg_nxt[4]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[4]~q ),
	.prn(vcc));
defparam \W_ipending_reg[4] .is_wysiwyg = "true";
defparam \W_ipending_reg[4] .power_up = "low";

cycloneive_lcell_comb \E_src1[3]~23 (
	.dataa(\D_iw[7]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[3]~23_combout ),
	.cout());
defparam \E_src1[3]~23 .lut_mask = 16'hAACC;
defparam \E_src1[3]~23 .sum_lutc_input = "datac";

dffeas \E_src1[3] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[3]~23_combout ),
	.asdata(\F_pc_plus_one[1]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

dffeas \W_ienable_reg[3] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~0_combout ),
	.q(\W_ienable_reg[3]~q ),
	.prn(vcc));
defparam \W_ienable_reg[3] .is_wysiwyg = "true";
defparam \W_ienable_reg[3] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[3]~1 (
	.dataa(\W_ienable_reg[3]~q ),
	.datab(dreg_1),
	.datac(gnd),
	.datad(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[3]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[3]~1_combout ),
	.cout());
defparam \W_ipending_reg_nxt[3]~1 .lut_mask = 16'hEEFF;
defparam \W_ipending_reg_nxt[3]~1 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[3] (
	.clk(wire_pll7_clk_0),
	.d(\W_ipending_reg_nxt[3]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[3]~q ),
	.prn(vcc));
defparam \W_ipending_reg[3] .is_wysiwyg = "true";
defparam \W_ipending_reg[3] .power_up = "low";

cycloneive_lcell_comb \E_src1[2]~24 (
	.dataa(\D_iw[6]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[2]~24_combout ),
	.cout());
defparam \E_src1[2]~24 .lut_mask = 16'hAACC;
defparam \E_src1[2]~24 .sum_lutc_input = "datac";

dffeas \E_src1[2] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[2]~24_combout ),
	.asdata(\F_pc_plus_one[0]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

dffeas \W_ienable_reg[2] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~0_combout ),
	.q(\W_ienable_reg[2]~q ),
	.prn(vcc));
defparam \W_ienable_reg[2] .is_wysiwyg = "true";
defparam \W_ienable_reg[2] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[2]~2 (
	.dataa(\W_ienable_reg[2]~q ),
	.datab(timeout_occurred),
	.datac(control_register_0),
	.datad(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[2]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[2]~2_combout ),
	.cout());
defparam \W_ipending_reg_nxt[2]~2 .lut_mask = 16'hFEFF;
defparam \W_ipending_reg_nxt[2]~2 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[2] (
	.clk(wire_pll7_clk_0),
	.d(\W_ipending_reg_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[2]~q ),
	.prn(vcc));
defparam \W_ipending_reg[2] .is_wysiwyg = "true";
defparam \W_ipending_reg[2] .power_up = "low";

cycloneive_lcell_comb \R_src1[1]~16 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\R_src1~15_combout ),
	.cin(gnd),
	.combout(\R_src1[1]~16_combout ),
	.cout());
defparam \R_src1[1]~16 .lut_mask = 16'hF7FF;
defparam \R_src1[1]~16 .sum_lutc_input = "datac";

dffeas \E_src1[1] (
	.clk(wire_pll7_clk_0),
	.d(\R_src1[1]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

dffeas \W_ienable_reg[1] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~0_combout ),
	.q(\W_ienable_reg[1]~q ),
	.prn(vcc));
defparam \W_ienable_reg[1] .is_wysiwyg = "true";
defparam \W_ienable_reg[1] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[1]~3 (
	.dataa(\W_ienable_reg[1]~q ),
	.datab(dreg_11),
	.datac(gnd),
	.datad(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[1]~3_combout ),
	.cout());
defparam \W_ipending_reg_nxt[1]~3 .lut_mask = 16'hEEFF;
defparam \W_ipending_reg_nxt[1]~3 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[1] (
	.clk(wire_pll7_clk_0),
	.d(\W_ipending_reg_nxt[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[1]~q ),
	.prn(vcc));
defparam \W_ipending_reg[1] .is_wysiwyg = "true";
defparam \W_ipending_reg[1] .power_up = "low";

cycloneive_lcell_comb \D_iw[1]~0 (
	.dataa(\W_ipending_reg[4]~q ),
	.datab(\W_ipending_reg[3]~q ),
	.datac(\W_ipending_reg[2]~q ),
	.datad(\W_ipending_reg[1]~q ),
	.cin(gnd),
	.combout(\D_iw[1]~0_combout ),
	.cout());
defparam \D_iw[1]~0 .lut_mask = 16'h7FFF;
defparam \D_iw[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[0]~17 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\R_src1~15_combout ),
	.cin(gnd),
	.combout(\R_src1[0]~17_combout ),
	.cout());
defparam \R_src1[0]~17 .lut_mask = 16'hF7FF;
defparam \R_src1[0]~17 .sum_lutc_input = "datac";

dffeas \E_src1[0] (
	.clk(wire_pll7_clk_0),
	.d(\R_src1[0]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

dffeas \W_ienable_reg[0] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~0_combout ),
	.q(\W_ienable_reg[0]~q ),
	.prn(vcc));
defparam \W_ienable_reg[0] .is_wysiwyg = "true";
defparam \W_ienable_reg[0] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[0]~4 (
	.dataa(\W_ienable_reg[0]~q ),
	.datab(irq1),
	.datac(gnd),
	.datad(\the_niosII_cpu_cpu_nios2_oci|the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[0]~4_combout ),
	.cout());
defparam \W_ipending_reg_nxt[0]~4 .lut_mask = 16'hEEFF;
defparam \W_ipending_reg_nxt[0]~4 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[0] (
	.clk(wire_pll7_clk_0),
	.d(\W_ipending_reg_nxt[0]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[0]~q ),
	.prn(vcc));
defparam \W_ipending_reg[0] .is_wysiwyg = "true";
defparam \W_ipending_reg[0] .power_up = "low";

cycloneive_lcell_comb \E_wrctl_estatus~0 (
	.dataa(\D_iw[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[7]~q ),
	.cin(gnd),
	.combout(\E_wrctl_estatus~0_combout ),
	.cout());
defparam \E_wrctl_estatus~0 .lut_mask = 16'hAAFF;
defparam \E_wrctl_estatus~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_wrctl_status~1 (
	.dataa(\R_ctrl_wrctl_inst~q ),
	.datab(\D_iw[9]~q ),
	.datac(\D_iw[10]~q ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\E_wrctl_status~1_combout ),
	.cout());
defparam \E_wrctl_status~1 .lut_mask = 16'hBFFF;
defparam \E_wrctl_status~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_estatus_reg_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_estatus_reg~q ),
	.datac(\E_wrctl_estatus~0_combout ),
	.datad(\E_wrctl_status~1_combout ),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~0 .lut_mask = 16'hEFFE;
defparam \W_estatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~7 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~7_combout ),
	.cout());
defparam \D_ctrl_exception~7 .lut_mask = 16'hEBBE;
defparam \D_ctrl_exception~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~24 (
	.dataa(\D_ctrl_exception~7_combout ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_exception~24_combout ),
	.cout());
defparam \D_ctrl_exception~24 .lut_mask = 16'hFEFE;
defparam \D_ctrl_exception~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~10 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~10_combout ),
	.cout());
defparam \D_ctrl_exception~10 .lut_mask = 16'hFBFF;
defparam \D_ctrl_exception~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~11 (
	.dataa(\D_iw[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~11_combout ),
	.cout());
defparam \D_ctrl_exception~11 .lut_mask = 16'hAAFF;
defparam \D_ctrl_exception~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~12 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_ctrl_exception~24_combout ),
	.datac(\D_ctrl_exception~10_combout ),
	.datad(\D_ctrl_exception~11_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~12_combout ),
	.cout());
defparam \D_ctrl_exception~12 .lut_mask = 16'hFFFE;
defparam \D_ctrl_exception~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~0 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~14_combout ),
	.datac(\Equal0~10_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_implicit_dst_eretaddr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~1 (
	.dataa(\Equal0~3_combout ),
	.datab(\Equal0~2_combout ),
	.datac(\Equal0~13_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~1 .lut_mask = 16'hBFFF;
defparam \D_ctrl_implicit_dst_eretaddr~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~2 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datab(\D_ctrl_force_src2_zero~0_combout ),
	.datac(\Equal0~14_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~2 .lut_mask = 16'hEFFF;
defparam \D_ctrl_implicit_dst_eretaddr~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~22 (
	.dataa(\D_ctrl_exception~12_combout ),
	.datab(\D_ctrl_exception~17_combout ),
	.datac(\D_ctrl_exception~21_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~22_combout ),
	.cout());
defparam \D_ctrl_exception~22 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~22 .sum_lutc_input = "datac";

dffeas R_ctrl_exception(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_exception~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_exception~q ),
	.prn(vcc));
defparam R_ctrl_exception.is_wysiwyg = "true";
defparam R_ctrl_exception.power_up = "low";

cycloneive_lcell_comb \W_estatus_reg_inst_nxt~1 (
	.dataa(\W_status_reg_pie~q ),
	.datab(\W_estatus_reg_inst_nxt~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~1 .lut_mask = 16'hAACC;
defparam \W_estatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

dffeas W_estatus_reg(
	.clk(wire_pll7_clk_0),
	.d(\W_estatus_reg_inst_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_estatus_reg~q ),
	.prn(vcc));
defparam W_estatus_reg.is_wysiwyg = "true";
defparam W_estatus_reg.power_up = "low";

cycloneive_lcell_comb \E_wrctl_bstatus~0 (
	.dataa(\D_iw[7]~q ),
	.datab(\E_wrctl_status~1_combout ),
	.datac(gnd),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_wrctl_bstatus~0_combout ),
	.cout());
defparam \E_wrctl_bstatus~0 .lut_mask = 16'hEEFF;
defparam \E_wrctl_bstatus~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_break~0 (
	.dataa(\D_iw[13]~q ),
	.datab(\D_iw[16]~q ),
	.datac(\D_op_opx_rsv17~0_combout ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.cout());
defparam \D_ctrl_break~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_break~0 .sum_lutc_input = "datac";

dffeas R_ctrl_break(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_break~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_break~q ),
	.prn(vcc));
defparam R_ctrl_break.is_wysiwyg = "true";
defparam R_ctrl_break.power_up = "low";

cycloneive_lcell_comb \W_bstatus_reg_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_bstatus_reg~q ),
	.datac(\E_wrctl_bstatus~0_combout ),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~0 .lut_mask = 16'hACFF;
defparam \W_bstatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_bstatus_reg_inst_nxt~1 (
	.dataa(\W_bstatus_reg_inst_nxt~0_combout ),
	.datab(\R_ctrl_break~q ),
	.datac(\W_status_reg_pie~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~1 .lut_mask = 16'hFEFE;
defparam \W_bstatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

dffeas W_bstatus_reg(
	.clk(wire_pll7_clk_0),
	.d(\W_bstatus_reg_inst_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_bstatus_reg~q ),
	.prn(vcc));
defparam W_bstatus_reg.is_wysiwyg = "true";
defparam W_bstatus_reg.power_up = "low";

cycloneive_lcell_comb \E_wrctl_status~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[7]~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_wrctl_status~0_combout ),
	.cout());
defparam \E_wrctl_status~0 .lut_mask = 16'h0FFF;
defparam \E_wrctl_status~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_status_reg_pie~q ),
	.datac(\E_wrctl_status~0_combout ),
	.datad(\E_wrctl_status~1_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~0_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~0 .lut_mask = 16'hEFFE;
defparam \W_status_reg_pie_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~1 (
	.dataa(\W_bstatus_reg~q ),
	.datab(\W_status_reg_pie_inst_nxt~0_combout ),
	.datac(\D_op_cmpge~0_combout ),
	.datad(\Equal62~9_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~1_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~1 .lut_mask = 16'hEFFE;
defparam \W_status_reg_pie_inst_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb D_op_eret(
	.dataa(\Equal0~8_combout ),
	.datab(\Equal62~9_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_eret~combout ),
	.cout());
defparam D_op_eret.lut_mask = 16'hEFFF;
defparam D_op_eret.sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_sel_nxt.10~0 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\R_ctrl_break~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_pc_sel_nxt.10~0_combout ),
	.cout());
defparam \F_pc_sel_nxt.10~0 .lut_mask = 16'hEEEE;
defparam \F_pc_sel_nxt.10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~2 (
	.dataa(\W_estatus_reg~q ),
	.datab(\W_status_reg_pie_inst_nxt~1_combout ),
	.datac(\D_op_eret~combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~2_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~2 .lut_mask = 16'hACFF;
defparam \W_status_reg_pie_inst_nxt~2 .sum_lutc_input = "datac";

dffeas W_status_reg_pie(
	.clk(wire_pll7_clk_0),
	.d(\W_status_reg_pie_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_status_reg_pie~q ),
	.prn(vcc));
defparam W_status_reg_pie.is_wysiwyg = "true";
defparam W_status_reg_pie.power_up = "low";

cycloneive_lcell_comb \D_iw[1]~1 (
	.dataa(\D_iw[1]~0_combout ),
	.datab(gnd),
	.datac(\W_ipending_reg[0]~q ),
	.datad(\W_status_reg_pie~q ),
	.cin(gnd),
	.combout(\D_iw[1]~1_combout ),
	.cout());
defparam \D_iw[1]~1 .lut_mask = 16'hAFFF;
defparam \D_iw[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_iw[1]~2 (
	.dataa(\D_iw[1]~1_combout ),
	.datab(hbreak_enabled1),
	.datac(gnd),
	.datad(\hbreak_req~0_combout ),
	.cin(gnd),
	.combout(\D_iw[1]~2_combout ),
	.cout());
defparam \D_iw[1]~2 .lut_mask = 16'hEEFF;
defparam \D_iw[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[11]~17 (
	.dataa(\F_iw[11]~16_combout ),
	.datab(src1_valid1),
	.datac(src_data_11),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[11]~17_combout ),
	.cout());
defparam \F_iw[11]~17 .lut_mask = 16'hFEFF;
defparam \F_iw[11]~17 .sum_lutc_input = "datac";

dffeas \D_iw[11] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[11]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

cycloneive_lcell_comb \Equal62~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~0_combout ),
	.cout());
defparam \Equal62~0 .lut_mask = 16'h7FFF;
defparam \Equal62~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~5 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'hFFBF;
defparam \Equal0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~8 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~5_combout ),
	.datad(\D_ctrl_alu_force_xor~14_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~8_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~8 .lut_mask = 16'h27FF;
defparam \D_ctrl_alu_subtract~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~9 (
	.dataa(\Equal62~0_combout ),
	.datab(\D_op_cmpge~0_combout ),
	.datac(gnd),
	.datad(\D_ctrl_alu_subtract~8_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~9_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~9 .lut_mask = 16'hEEFF;
defparam \D_ctrl_alu_subtract~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~5 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\D_iw[11]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~5_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~5 .lut_mask = 16'hFF96;
defparam \D_ctrl_alu_subtract~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~10 (
	.dataa(\D_ctrl_alu_subtract~5_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~10_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~10 .lut_mask = 16'hBFBF;
defparam \D_ctrl_alu_subtract~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_alu_sub~0 (
	.dataa(\R_valid~q ),
	.datab(\D_ctrl_alu_subtract~9_combout ),
	.datac(\Equal0~8_combout ),
	.datad(\D_ctrl_alu_subtract~10_combout ),
	.cin(gnd),
	.combout(\E_alu_sub~0_combout ),
	.cout());
defparam \E_alu_sub~0 .lut_mask = 16'hFFFE;
defparam \E_alu_sub~0 .sum_lutc_input = "datac";

dffeas E_alu_sub(
	.clk(wire_pll7_clk_0),
	.d(\E_alu_sub~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_alu_sub~q ),
	.prn(vcc));
defparam E_alu_sub.is_wysiwyg = "true";
defparam E_alu_sub.power_up = "low";

cycloneive_lcell_comb \E_src2[5]~15 (
	.dataa(\R_ctrl_src_imm5_shift_rot~q ),
	.datab(\R_ctrl_hi_imm16~q ),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_src2[5]~15_combout ),
	.cout());
defparam \E_src2[5]~15 .lut_mask = 16'hFEFE;
defparam \E_src2[5]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[6]~0 (
	.dataa(\D_iw[12]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[6]~0_combout ),
	.cout());
defparam \R_src2_lo[6]~0 .lut_mask = 16'hACFF;
defparam \R_src2_lo[6]~0 .sum_lutc_input = "datac";

dffeas \E_src2[6] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[6]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[6]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[6]~20 (
	.dataa(\D_iw[10]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[6]~20_combout ),
	.cout());
defparam \E_src1[6]~20 .lut_mask = 16'hAACC;
defparam \E_src1[6]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[3]~6 (
	.dataa(F_pc_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[2]~5 ),
	.combout(\F_pc_plus_one[3]~6_combout ),
	.cout(\F_pc_plus_one[3]~7 ));
defparam \F_pc_plus_one[3]~6 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[4]~8 (
	.dataa(F_pc_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[3]~7 ),
	.combout(\F_pc_plus_one[4]~8_combout ),
	.cout(\F_pc_plus_one[4]~9 ));
defparam \F_pc_plus_one[4]~8 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[4]~8 .sum_lutc_input = "cin";

dffeas \E_src1[6] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[6]~20_combout ),
	.asdata(\F_pc_plus_one[4]~8_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[5]~1 (
	.dataa(\D_iw[11]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[5]~1_combout ),
	.cout());
defparam \R_src2_lo[5]~1 .lut_mask = 16'hACFF;
defparam \R_src2_lo[5]~1 .sum_lutc_input = "datac";

dffeas \E_src2[5] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[5]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_src2[5]~q ),
	.datad(\E_alu_sub~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h0FF0;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[5]~21 (
	.dataa(\D_iw[9]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[5]~21_combout ),
	.cout());
defparam \E_src1[5]~21 .lut_mask = 16'hAACC;
defparam \E_src1[5]~21 .sum_lutc_input = "datac";

dffeas \E_src1[5] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[5]~21_combout ),
	.asdata(\F_pc_plus_one[3]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[4]~q ),
	.cin(gnd),
	.combout(\Add1~2_combout ),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[3]~q ),
	.cin(gnd),
	.combout(\Add1~3_combout ),
	.cout());
defparam \Add1~3 .lut_mask = 16'h0FF0;
defparam \Add1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[2]~q ),
	.cin(gnd),
	.combout(\Add1~4_combout ),
	.cout());
defparam \Add1~4 .lut_mask = 16'h0FF0;
defparam \Add1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[1]~q ),
	.cin(gnd),
	.combout(\Add1~5_combout ),
	.cout());
defparam \Add1~5 .lut_mask = 16'h0FF0;
defparam \Add1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[0]~q ),
	.cin(gnd),
	.combout(\Add1~6_combout ),
	.cout());
defparam \Add1~6 .lut_mask = 16'h0FF0;
defparam \Add1~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~8 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add1~8_cout ));
defparam \Add1~8 .lut_mask = 16'h00AA;
defparam \Add1~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~9 (
	.dataa(\Add1~6_combout ),
	.datab(\E_src1[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~8_cout ),
	.combout(\Add1~9_combout ),
	.cout(\Add1~10 ));
defparam \Add1~9 .lut_mask = 16'h967F;
defparam \Add1~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~11 (
	.dataa(\Add1~5_combout ),
	.datab(\E_src1[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~10 ),
	.combout(\Add1~11_combout ),
	.cout(\Add1~12 ));
defparam \Add1~11 .lut_mask = 16'h96EF;
defparam \Add1~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~13 (
	.dataa(\Add1~4_combout ),
	.datab(\E_src1[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~12 ),
	.combout(\Add1~13_combout ),
	.cout(\Add1~14 ));
defparam \Add1~13 .lut_mask = 16'h967F;
defparam \Add1~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~15 (
	.dataa(\Add1~3_combout ),
	.datab(\E_src1[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~14 ),
	.combout(\Add1~15_combout ),
	.cout(\Add1~16 ));
defparam \Add1~15 .lut_mask = 16'h96EF;
defparam \Add1~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~17 (
	.dataa(\Add1~2_combout ),
	.datab(\E_src1[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~16 ),
	.combout(\Add1~17_combout ),
	.cout(\Add1~18 ));
defparam \Add1~17 .lut_mask = 16'h967F;
defparam \Add1~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~19 (
	.dataa(\Add1~1_combout ),
	.datab(\E_src1[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~18 ),
	.combout(\Add1~19_combout ),
	.cout(\Add1~20 ));
defparam \Add1~19 .lut_mask = 16'h96EF;
defparam \Add1~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~21 (
	.dataa(\Add1~0_combout ),
	.datab(\E_src1[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~20 ),
	.combout(\Add1~21_combout ),
	.cout(\Add1~22 ));
defparam \Add1~21 .lut_mask = 16'h967F;
defparam \Add1~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \D_logic_op_raw[1]~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_logic_op_raw[1]~0_combout ),
	.cout());
defparam \D_logic_op_raw[1]~0 .lut_mask = 16'hEFFF;
defparam \D_logic_op_raw[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~10 (
	.dataa(\Equal62~0_combout ),
	.datab(\D_op_cmpge~0_combout ),
	.datac(\D_ctrl_alu_force_xor~14_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~10_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~10 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~11 (
	.dataa(\Equal0~5_combout ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~4_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~11_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~11 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~13 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~13_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~13 .lut_mask = 16'hFFD8;
defparam \D_ctrl_alu_force_xor~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~12 (
	.dataa(\D_ctrl_alu_force_xor~10_combout ),
	.datab(\D_ctrl_alu_force_xor~11_combout ),
	.datac(\Equal0~8_combout ),
	.datad(\D_ctrl_alu_force_xor~13_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~12_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~12 .lut_mask = 16'hFFFE;
defparam \D_ctrl_alu_force_xor~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_logic_op[1]~0 (
	.dataa(\D_logic_op_raw[1]~0_combout ),
	.datab(\D_ctrl_alu_force_xor~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.cout());
defparam \D_logic_op[1]~0 .lut_mask = 16'hEEEE;
defparam \D_logic_op[1]~0 .sum_lutc_input = "datac";

dffeas \R_logic_op[1] (
	.clk(wire_pll7_clk_0),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[1]~q ),
	.prn(vcc));
defparam \R_logic_op[1] .is_wysiwyg = "true";
defparam \R_logic_op[1] .power_up = "low";

cycloneive_lcell_comb \D_logic_op[0]~1 (
	.dataa(\D_ctrl_alu_force_xor~12_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\Equal0~8_combout ),
	.cin(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.cout());
defparam \D_logic_op[0]~1 .lut_mask = 16'hFAFC;
defparam \D_logic_op[0]~1 .sum_lutc_input = "datac";

dffeas \R_logic_op[0] (
	.clk(wire_pll7_clk_0),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[0]~q ),
	.prn(vcc));
defparam \R_logic_op[0] .is_wysiwyg = "true";
defparam \R_logic_op[0] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[6]~0 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[6]~q ),
	.datac(\E_src1[6]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[6]~0_combout ),
	.cout());
defparam \E_logic_result[6]~0 .lut_mask = 16'h6996;
defparam \E_logic_result[6]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~9 (
	.dataa(\D_iw[13]~q ),
	.datab(gnd),
	.datac(\D_iw[11]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
defparam \Equal0~9 .lut_mask = 16'hAFFF;
defparam \Equal0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~11 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~11_combout ),
	.cout());
defparam \Equal0~11 .lut_mask = 16'hFFF7;
defparam \Equal0~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_logic~0 (
	.dataa(gnd),
	.datab(\D_iw[4]~q ),
	.datac(\Equal0~10_combout ),
	.datad(\Equal0~11_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.cout());
defparam \D_ctrl_logic~0 .lut_mask = 16'h3FFF;
defparam \D_ctrl_logic~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb D_ctrl_logic(
	.dataa(\Equal0~8_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\Equal0~9_combout ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~combout ),
	.cout());
defparam D_ctrl_logic.lut_mask = 16'hFEFF;
defparam D_ctrl_logic.sum_lutc_input = "datac";

dffeas R_ctrl_logic(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_logic~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_logic~q ),
	.prn(vcc));
defparam R_ctrl_logic.is_wysiwyg = "true";
defparam R_ctrl_logic.power_up = "low";

cycloneive_lcell_comb \W_alu_result[6]~20 (
	.dataa(\Add1~21_combout ),
	.datab(\E_logic_result[6]~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[6]~20_combout ),
	.cout());
defparam \W_alu_result[6]~20 .lut_mask = 16'hAACC;
defparam \W_alu_result[6]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot_right~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot_right~1 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_shift_rot_right~0_combout ),
	.datad(\D_iw[13]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~1 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot_right(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_shift_rot_right~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam R_ctrl_shift_rot_right.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[5]~18 (
	.dataa(\E_shift_rot_result[6]~q ),
	.datab(\E_shift_rot_result[4]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[5]~18_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[5]~18 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[5]~18 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[5] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[5]~18_combout ),
	.asdata(\E_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[5] .is_wysiwyg = "true";
defparam \E_shift_rot_result[5] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[4]~22 (
	.dataa(\E_shift_rot_result[5]~q ),
	.datab(\E_shift_rot_result[3]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[4]~22_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[4]~22 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[4]~22 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[4] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[4]~22_combout ),
	.asdata(\E_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[4] .is_wysiwyg = "true";
defparam \E_shift_rot_result[4] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[3]~23 (
	.dataa(\E_shift_rot_result[4]~q ),
	.datab(\E_shift_rot_result[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[3]~23_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[3]~23 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[3]~23 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[3] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[3]~23_combout ),
	.asdata(\E_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[3] .is_wysiwyg = "true";
defparam \E_shift_rot_result[3] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[2]~24 (
	.dataa(\E_shift_rot_result[3]~q ),
	.datab(\E_shift_rot_result[1]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[2]~24_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[2]~24 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[2]~24 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[2] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[2]~24_combout ),
	.asdata(\E_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[2] .is_wysiwyg = "true";
defparam \E_shift_rot_result[2] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[1]~26 (
	.dataa(\E_shift_rot_result[2]~q ),
	.datab(\E_shift_rot_result[0]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[1]~26_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[1]~26 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[1]~26 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[1] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[1]~26_combout ),
	.asdata(\E_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[1] .is_wysiwyg = "true";
defparam \E_shift_rot_result[1] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[0]~28 (
	.dataa(\E_shift_rot_result[1]~q ),
	.datab(\E_shift_rot_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[0]~28_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[0]~28 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[0]~28 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[0] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[0]~28_combout ),
	.asdata(\E_src1[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[0] .is_wysiwyg = "true";
defparam \E_shift_rot_result[0] .power_up = "low";

cycloneive_lcell_comb \R_ctrl_rot_right_nxt~0 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~7_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\R_ctrl_rot_right_nxt~0_combout ),
	.cout());
defparam \R_ctrl_rot_right_nxt~0 .lut_mask = 16'hFEFF;
defparam \R_ctrl_rot_right_nxt~0 .sum_lutc_input = "datac";

dffeas R_ctrl_rot_right(
	.clk(wire_pll7_clk_0),
	.d(\R_ctrl_rot_right_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_rot_right.is_wysiwyg = "true";
defparam R_ctrl_rot_right.power_up = "low";

cycloneive_lcell_comb \D_ctrl_shift_logical~1 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~4_combout ),
	.datad(\Equal62~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~1_combout ),
	.cout());
defparam \D_ctrl_shift_logical~1 .lut_mask = 16'hFFB8;
defparam \D_ctrl_shift_logical~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_logical~2 (
	.dataa(\Equal0~8_combout ),
	.datab(\D_iw[15]~q ),
	.datac(\D_ctrl_shift_logical~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~2_combout ),
	.cout());
defparam \D_ctrl_shift_logical~2 .lut_mask = 16'hFEFE;
defparam \D_ctrl_shift_logical~2 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_logical(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_shift_logical~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_logical~q ),
	.prn(vcc));
defparam R_ctrl_shift_logical.is_wysiwyg = "true";
defparam R_ctrl_shift_logical.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_fill_bit~0 (
	.dataa(\E_shift_rot_result[0]~q ),
	.datab(\E_shift_rot_result[31]~q ),
	.datac(\R_ctrl_rot_right~q ),
	.datad(\R_ctrl_shift_logical~q ),
	.cin(gnd),
	.combout(\E_shift_rot_fill_bit~0_combout ),
	.cout());
defparam \E_shift_rot_fill_bit~0 .lut_mask = 16'hACFF;
defparam \E_shift_rot_fill_bit~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_shift_rot_result_nxt[31]~30 (
	.dataa(\E_shift_rot_fill_bit~0_combout ),
	.datab(\E_shift_rot_result[30]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[31]~30_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[31]~30 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[31]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[31]~18 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.datad(\R_src1~15_combout ),
	.cin(gnd),
	.combout(\R_src1[31]~18_combout ),
	.cout());
defparam \R_src1[31]~18 .lut_mask = 16'hF7FF;
defparam \R_src1[31]~18 .sum_lutc_input = "datac";

dffeas \E_src1[31] (
	.clk(wire_pll7_clk_0),
	.d(\R_src1[31]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

dffeas \E_shift_rot_result[31] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[31]~30_combout ),
	.asdata(\E_src1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[31] .is_wysiwyg = "true";
defparam \E_shift_rot_result[31] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[30]~31 (
	.dataa(\E_shift_rot_result[31]~q ),
	.datab(\E_shift_rot_result[29]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[30]~31_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[30]~31 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[30]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[30]~19 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.datad(\R_src1~15_combout ),
	.cin(gnd),
	.combout(\R_src1[30]~19_combout ),
	.cout());
defparam \R_src1[30]~19 .lut_mask = 16'hF7FF;
defparam \R_src1[30]~19 .sum_lutc_input = "datac";

dffeas \E_src1[30] (
	.clk(wire_pll7_clk_0),
	.d(\R_src1[30]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

dffeas \E_shift_rot_result[30] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[30]~31_combout ),
	.asdata(\E_src1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[30] .is_wysiwyg = "true";
defparam \E_shift_rot_result[30] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[29]~29 (
	.dataa(\E_shift_rot_result[30]~q ),
	.datab(\E_shift_rot_result[28]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[29]~29_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[29]~29 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[29]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[29]~20 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.datad(\R_src1~15_combout ),
	.cin(gnd),
	.combout(\R_src1[29]~20_combout ),
	.cout());
defparam \R_src1[29]~20 .lut_mask = 16'hF7FF;
defparam \R_src1[29]~20 .sum_lutc_input = "datac";

dffeas \E_src1[29] (
	.clk(wire_pll7_clk_0),
	.d(\R_src1[29]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

dffeas \E_shift_rot_result[29] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[29]~29_combout ),
	.asdata(\E_src1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[29] .is_wysiwyg = "true";
defparam \E_shift_rot_result[29] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[28]~27 (
	.dataa(\E_shift_rot_result[29]~q ),
	.datab(\E_shift_rot_result[27]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[28]~27_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[28]~27 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[28]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[28]~21 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.datad(\R_src1~15_combout ),
	.cin(gnd),
	.combout(\R_src1[28]~21_combout ),
	.cout());
defparam \R_src1[28]~21 .lut_mask = 16'hF7FF;
defparam \R_src1[28]~21 .sum_lutc_input = "datac";

dffeas \E_src1[28] (
	.clk(wire_pll7_clk_0),
	.d(\R_src1[28]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

dffeas \E_shift_rot_result[28] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[28]~27_combout ),
	.asdata(\E_src1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[28] .is_wysiwyg = "true";
defparam \E_shift_rot_result[28] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[27]~25 (
	.dataa(\E_shift_rot_result[28]~q ),
	.datab(\E_shift_rot_result[26]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[27]~25_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[27]~25 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[27]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[27]~22 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.datad(\R_src1~15_combout ),
	.cin(gnd),
	.combout(\R_src1[27]~22_combout ),
	.cout());
defparam \R_src1[27]~22 .lut_mask = 16'hF7FF;
defparam \R_src1[27]~22 .sum_lutc_input = "datac";

dffeas \E_src1[27] (
	.clk(wire_pll7_clk_0),
	.d(\R_src1[27]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

dffeas \E_shift_rot_result[27] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[27]~25_combout ),
	.asdata(\E_src1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[27] .is_wysiwyg = "true";
defparam \E_shift_rot_result[27] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[26]~1 (
	.dataa(\E_shift_rot_result[27]~q ),
	.datab(\E_shift_rot_result[25]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[26]~1_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[26]~1 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[26]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[30]~49 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_30),
	.datad(out_data_buffer_30),
	.cin(gnd),
	.combout(\F_iw[30]~49_combout ),
	.cout());
defparam \F_iw[30]~49 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[30]~50 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[30]~49_combout ),
	.datac(src_payload),
	.datad(out_payload_14),
	.cin(gnd),
	.combout(\F_iw[30]~50_combout ),
	.cout());
defparam \F_iw[30]~50 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~50 .sum_lutc_input = "datac";

dffeas \D_iw[30] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[30]~50_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

cycloneive_lcell_comb \E_src1[26]~0 (
	.dataa(\D_iw[30]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[26]~0_combout ),
	.cout());
defparam \E_src1[26]~0 .lut_mask = 16'hAACC;
defparam \E_src1[26]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[5]~10 (
	.dataa(F_pc_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[4]~9 ),
	.combout(\F_pc_plus_one[5]~10_combout ),
	.cout(\F_pc_plus_one[5]~11 ));
defparam \F_pc_plus_one[5]~10 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[5]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[6]~12 (
	.dataa(F_pc_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[5]~11 ),
	.combout(\F_pc_plus_one[6]~12_combout ),
	.cout(\F_pc_plus_one[6]~13 ));
defparam \F_pc_plus_one[6]~12 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[6]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[7]~14 (
	.dataa(F_pc_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[6]~13 ),
	.combout(\F_pc_plus_one[7]~14_combout ),
	.cout(\F_pc_plus_one[7]~15 ));
defparam \F_pc_plus_one[7]~14 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[7]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[8]~16 (
	.dataa(F_pc_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[7]~15 ),
	.combout(\F_pc_plus_one[8]~16_combout ),
	.cout(\F_pc_plus_one[8]~17 ));
defparam \F_pc_plus_one[8]~16 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[8]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[9]~18 (
	.dataa(F_pc_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[8]~17 ),
	.combout(\F_pc_plus_one[9]~18_combout ),
	.cout(\F_pc_plus_one[9]~19 ));
defparam \F_pc_plus_one[9]~18 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[9]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[10]~20 (
	.dataa(F_pc_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[9]~19 ),
	.combout(\F_pc_plus_one[10]~20_combout ),
	.cout(\F_pc_plus_one[10]~21 ));
defparam \F_pc_plus_one[10]~20 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[10]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[11]~22 (
	.dataa(F_pc_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[10]~21 ),
	.combout(\F_pc_plus_one[11]~22_combout ),
	.cout(\F_pc_plus_one[11]~23 ));
defparam \F_pc_plus_one[11]~22 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[11]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[12]~24 (
	.dataa(F_pc_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[11]~23 ),
	.combout(\F_pc_plus_one[12]~24_combout ),
	.cout(\F_pc_plus_one[12]~25 ));
defparam \F_pc_plus_one[12]~24 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[12]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[13]~26 (
	.dataa(F_pc_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[12]~25 ),
	.combout(\F_pc_plus_one[13]~26_combout ),
	.cout(\F_pc_plus_one[13]~27 ));
defparam \F_pc_plus_one[13]~26 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[13]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[14]~28 (
	.dataa(F_pc_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[13]~27 ),
	.combout(\F_pc_plus_one[14]~28_combout ),
	.cout(\F_pc_plus_one[14]~29 ));
defparam \F_pc_plus_one[14]~28 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[14]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[15]~30 (
	.dataa(F_pc_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[14]~29 ),
	.combout(\F_pc_plus_one[15]~30_combout ),
	.cout(\F_pc_plus_one[15]~31 ));
defparam \F_pc_plus_one[15]~30 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[15]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[16]~32 (
	.dataa(F_pc_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[15]~31 ),
	.combout(\F_pc_plus_one[16]~32_combout ),
	.cout(\F_pc_plus_one[16]~33 ));
defparam \F_pc_plus_one[16]~32 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[16]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[17]~34 (
	.dataa(F_pc_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[16]~33 ),
	.combout(\F_pc_plus_one[17]~34_combout ),
	.cout(\F_pc_plus_one[17]~35 ));
defparam \F_pc_plus_one[17]~34 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[17]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[18]~36 (
	.dataa(F_pc_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[17]~35 ),
	.combout(\F_pc_plus_one[18]~36_combout ),
	.cout(\F_pc_plus_one[18]~37 ));
defparam \F_pc_plus_one[18]~36 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[18]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[19]~38 (
	.dataa(F_pc_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[18]~37 ),
	.combout(\F_pc_plus_one[19]~38_combout ),
	.cout(\F_pc_plus_one[19]~39 ));
defparam \F_pc_plus_one[19]~38 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[19]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[20]~40 (
	.dataa(F_pc_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[19]~39 ),
	.combout(\F_pc_plus_one[20]~40_combout ),
	.cout(\F_pc_plus_one[20]~41 ));
defparam \F_pc_plus_one[20]~40 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[20]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[21]~42 (
	.dataa(F_pc_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[20]~41 ),
	.combout(\F_pc_plus_one[21]~42_combout ),
	.cout(\F_pc_plus_one[21]~43 ));
defparam \F_pc_plus_one[21]~42 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[21]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[22]~44 (
	.dataa(F_pc_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[21]~43 ),
	.combout(\F_pc_plus_one[22]~44_combout ),
	.cout(\F_pc_plus_one[22]~45 ));
defparam \F_pc_plus_one[22]~44 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[22]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[23]~46 (
	.dataa(F_pc_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[22]~45 ),
	.combout(\F_pc_plus_one[23]~46_combout ),
	.cout(\F_pc_plus_one[23]~47 ));
defparam \F_pc_plus_one[23]~46 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[23]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[24]~48 (
	.dataa(F_pc_24),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\F_pc_plus_one[23]~47 ),
	.combout(\F_pc_plus_one[24]~48_combout ),
	.cout());
defparam \F_pc_plus_one[24]~48 .lut_mask = 16'h5A5A;
defparam \F_pc_plus_one[24]~48 .sum_lutc_input = "cin";

dffeas \E_src1[26] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[26]~0_combout ),
	.asdata(\F_pc_plus_one[24]~48_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

dffeas \E_shift_rot_result[26] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[26]~1_combout ),
	.asdata(\E_src1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[26] .is_wysiwyg = "true";
defparam \E_shift_rot_result[26] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[25]~2 (
	.dataa(\E_shift_rot_result[26]~q ),
	.datab(\E_shift_rot_result[24]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[25]~2_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[25]~2 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[25]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[29]~51 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_29),
	.datad(out_data_buffer_29),
	.cin(gnd),
	.combout(\F_iw[29]~51_combout ),
	.cout());
defparam \F_iw[29]~51 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[29]~52 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[29]~51_combout ),
	.datac(out_payload_13),
	.datad(src_payload),
	.cin(gnd),
	.combout(\F_iw[29]~52_combout ),
	.cout());
defparam \F_iw[29]~52 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~52 .sum_lutc_input = "datac";

dffeas \D_iw[29] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[29]~52_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

cycloneive_lcell_comb \E_src1[25]~1 (
	.dataa(\D_iw[29]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[25]~1_combout ),
	.cout());
defparam \E_src1[25]~1 .lut_mask = 16'hAACC;
defparam \E_src1[25]~1 .sum_lutc_input = "datac";

dffeas \E_src1[25] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[25]~1_combout ),
	.asdata(\F_pc_plus_one[23]~46_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

dffeas \E_shift_rot_result[25] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[25]~2_combout ),
	.asdata(\E_src1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[25] .is_wysiwyg = "true";
defparam \E_shift_rot_result[25] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[24]~3 (
	.dataa(\E_shift_rot_result[25]~q ),
	.datab(\E_shift_rot_result[23]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[24]~3_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[24]~3 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[24]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[28]~53 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_28),
	.datad(out_data_buffer_28),
	.cin(gnd),
	.combout(\F_iw[28]~53_combout ),
	.cout());
defparam \F_iw[28]~53 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[28]~54 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[28]~53_combout ),
	.datac(src_payload),
	.datad(out_payload_12),
	.cin(gnd),
	.combout(\F_iw[28]~54_combout ),
	.cout());
defparam \F_iw[28]~54 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~54 .sum_lutc_input = "datac";

dffeas \D_iw[28] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[28]~54_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

cycloneive_lcell_comb \E_src1[24]~2 (
	.dataa(\D_iw[28]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[24]~2_combout ),
	.cout());
defparam \E_src1[24]~2 .lut_mask = 16'hAACC;
defparam \E_src1[24]~2 .sum_lutc_input = "datac";

dffeas \E_src1[24] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[24]~2_combout ),
	.asdata(\F_pc_plus_one[22]~44_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

dffeas \E_shift_rot_result[24] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[24]~3_combout ),
	.asdata(\E_src1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[24] .is_wysiwyg = "true";
defparam \E_shift_rot_result[24] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[23]~4 (
	.dataa(\E_shift_rot_result[24]~q ),
	.datab(\E_shift_rot_result[22]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[23]~4_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[23]~4 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[23]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[27]~55 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_27),
	.datad(out_data_buffer_27),
	.cin(gnd),
	.combout(\F_iw[27]~55_combout ),
	.cout());
defparam \F_iw[27]~55 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[27]~56 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[27]~55_combout ),
	.datac(out_payload_11),
	.datad(src_payload),
	.cin(gnd),
	.combout(\F_iw[27]~56_combout ),
	.cout());
defparam \F_iw[27]~56 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~56 .sum_lutc_input = "datac";

dffeas \D_iw[27] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[27]~56_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

cycloneive_lcell_comb \E_src1[23]~3 (
	.dataa(\D_iw[27]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[23]~3_combout ),
	.cout());
defparam \E_src1[23]~3 .lut_mask = 16'hAACC;
defparam \E_src1[23]~3 .sum_lutc_input = "datac";

dffeas \E_src1[23] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[23]~3_combout ),
	.asdata(\F_pc_plus_one[21]~42_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

dffeas \E_shift_rot_result[23] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[23]~4_combout ),
	.asdata(\E_src1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[23] .is_wysiwyg = "true";
defparam \E_shift_rot_result[23] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[22]~5 (
	.dataa(\E_shift_rot_result[23]~q ),
	.datab(\E_shift_rot_result[21]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[22]~5_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[22]~5 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[22]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[26]~57 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_26),
	.datad(out_data_buffer_26),
	.cin(gnd),
	.combout(\F_iw[26]~57_combout ),
	.cout());
defparam \F_iw[26]~57 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[26]~58 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[26]~57_combout ),
	.datac(src_payload),
	.datad(out_payload_10),
	.cin(gnd),
	.combout(\F_iw[26]~58_combout ),
	.cout());
defparam \F_iw[26]~58 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~58 .sum_lutc_input = "datac";

dffeas \D_iw[26] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[26]~58_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

cycloneive_lcell_comb \E_src1[22]~4 (
	.dataa(\D_iw[26]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[22]~4_combout ),
	.cout());
defparam \E_src1[22]~4 .lut_mask = 16'hAACC;
defparam \E_src1[22]~4 .sum_lutc_input = "datac";

dffeas \E_src1[22] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[22]~4_combout ),
	.asdata(\F_pc_plus_one[20]~40_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

dffeas \E_shift_rot_result[22] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[22]~5_combout ),
	.asdata(\E_src1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[22] .is_wysiwyg = "true";
defparam \E_shift_rot_result[22] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[21]~6 (
	.dataa(\E_shift_rot_result[22]~q ),
	.datab(\E_shift_rot_result[20]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[21]~6_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[21]~6 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[21]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[25]~59 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_25),
	.datad(out_data_buffer_25),
	.cin(gnd),
	.combout(\F_iw[25]~59_combout ),
	.cout());
defparam \F_iw[25]~59 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[25]~60 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[25]~59_combout ),
	.datac(src_payload),
	.datad(out_payload_9),
	.cin(gnd),
	.combout(\F_iw[25]~60_combout ),
	.cout());
defparam \F_iw[25]~60 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~60 .sum_lutc_input = "datac";

dffeas \D_iw[25] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[25]~60_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

cycloneive_lcell_comb \E_src1[21]~5 (
	.dataa(\D_iw[25]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[21]~5_combout ),
	.cout());
defparam \E_src1[21]~5 .lut_mask = 16'hAACC;
defparam \E_src1[21]~5 .sum_lutc_input = "datac";

dffeas \E_src1[21] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[21]~5_combout ),
	.asdata(\F_pc_plus_one[19]~38_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

dffeas \E_shift_rot_result[21] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[21]~6_combout ),
	.asdata(\E_src1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[21] .is_wysiwyg = "true";
defparam \E_shift_rot_result[21] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[20]~7 (
	.dataa(\E_shift_rot_result[21]~q ),
	.datab(\E_shift_rot_result[19]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[20]~7_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[20]~7 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[20]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[24]~61 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_24),
	.datad(out_data_buffer_24),
	.cin(gnd),
	.combout(\F_iw[24]~61_combout ),
	.cout());
defparam \F_iw[24]~61 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[24]~62 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[24]~61_combout ),
	.datac(src_payload),
	.datad(out_payload_8),
	.cin(gnd),
	.combout(\F_iw[24]~62_combout ),
	.cout());
defparam \F_iw[24]~62 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~62 .sum_lutc_input = "datac";

dffeas \D_iw[24] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[24]~62_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

cycloneive_lcell_comb \E_src1[20]~6 (
	.dataa(\D_iw[24]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[20]~6_combout ),
	.cout());
defparam \E_src1[20]~6 .lut_mask = 16'hAACC;
defparam \E_src1[20]~6 .sum_lutc_input = "datac";

dffeas \E_src1[20] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[20]~6_combout ),
	.asdata(\F_pc_plus_one[18]~36_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

dffeas \E_shift_rot_result[20] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[20]~7_combout ),
	.asdata(\E_src1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[20] .is_wysiwyg = "true";
defparam \E_shift_rot_result[20] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[19]~8 (
	.dataa(\E_shift_rot_result[20]~q ),
	.datab(\E_shift_rot_result[18]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[19]~8_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[19]~8 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[19]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[23]~63 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_23),
	.datad(out_data_buffer_23),
	.cin(gnd),
	.combout(\F_iw[23]~63_combout ),
	.cout());
defparam \F_iw[23]~63 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[23]~64 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[23]~63_combout ),
	.datac(src_payload),
	.datad(out_payload_7),
	.cin(gnd),
	.combout(\F_iw[23]~64_combout ),
	.cout());
defparam \F_iw[23]~64 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~64 .sum_lutc_input = "datac";

dffeas \D_iw[23] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[23]~64_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

cycloneive_lcell_comb \E_src1[19]~7 (
	.dataa(\D_iw[23]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[19]~7_combout ),
	.cout());
defparam \E_src1[19]~7 .lut_mask = 16'hAACC;
defparam \E_src1[19]~7 .sum_lutc_input = "datac";

dffeas \E_src1[19] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[19]~7_combout ),
	.asdata(\F_pc_plus_one[17]~34_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

dffeas \E_shift_rot_result[19] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[19]~8_combout ),
	.asdata(\E_src1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[19] .is_wysiwyg = "true";
defparam \E_shift_rot_result[19] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[18]~9 (
	.dataa(\E_shift_rot_result[19]~q ),
	.datab(\E_shift_rot_result[17]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[18]~9_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[18]~9 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[18]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[22]~65 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_22),
	.datad(out_data_buffer_22),
	.cin(gnd),
	.combout(\F_iw[22]~65_combout ),
	.cout());
defparam \F_iw[22]~65 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[22]~66 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[22]~65_combout ),
	.datac(src_payload),
	.datad(out_payload_6),
	.cin(gnd),
	.combout(\F_iw[22]~66_combout ),
	.cout());
defparam \F_iw[22]~66 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~66 .sum_lutc_input = "datac";

dffeas \D_iw[22] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[22]~66_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

cycloneive_lcell_comb \E_src1[18]~8 (
	.dataa(\D_iw[22]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[18]~8_combout ),
	.cout());
defparam \E_src1[18]~8 .lut_mask = 16'hAACC;
defparam \E_src1[18]~8 .sum_lutc_input = "datac";

dffeas \E_src1[18] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[18]~8_combout ),
	.asdata(\F_pc_plus_one[16]~32_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

dffeas \E_shift_rot_result[18] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[18]~9_combout ),
	.asdata(\E_src1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[18] .is_wysiwyg = "true";
defparam \E_shift_rot_result[18] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[17]~10 (
	.dataa(\E_shift_rot_result[18]~q ),
	.datab(\E_shift_rot_result[16]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[17]~10_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[17]~10 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[17]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[21]~47 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_21),
	.datad(out_data_buffer_21),
	.cin(gnd),
	.combout(\F_iw[21]~47_combout ),
	.cout());
defparam \F_iw[21]~47 .lut_mask = 16'hFFFE;
defparam \F_iw[21]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[21]~48 (
	.dataa(\F_iw[21]~47_combout ),
	.datab(out_payload_5),
	.datac(src_payload),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[21]~48_combout ),
	.cout());
defparam \F_iw[21]~48 .lut_mask = 16'hFEFF;
defparam \F_iw[21]~48 .sum_lutc_input = "datac";

dffeas \D_iw[21] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[21]~48_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cycloneive_lcell_comb \E_src1[17]~9 (
	.dataa(\D_iw[21]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[17]~9_combout ),
	.cout());
defparam \E_src1[17]~9 .lut_mask = 16'hAACC;
defparam \E_src1[17]~9 .sum_lutc_input = "datac";

dffeas \E_src1[17] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[17]~9_combout ),
	.asdata(\F_pc_plus_one[15]~30_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

dffeas \E_shift_rot_result[17] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[17]~10_combout ),
	.asdata(\E_src1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[17] .is_wysiwyg = "true";
defparam \E_shift_rot_result[17] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[16]~11 (
	.dataa(\E_shift_rot_result[17]~q ),
	.datab(\E_shift_rot_result[15]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[16]~11_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[16]~11 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[16]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[20]~67 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_20),
	.datad(out_data_buffer_20),
	.cin(gnd),
	.combout(\F_iw[20]~67_combout ),
	.cout());
defparam \F_iw[20]~67 .lut_mask = 16'hFFFE;
defparam \F_iw[20]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[20]~68 (
	.dataa(\F_iw[20]~67_combout ),
	.datab(out_payload_4),
	.datac(src_payload),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[20]~68_combout ),
	.cout());
defparam \F_iw[20]~68 .lut_mask = 16'hFEFF;
defparam \F_iw[20]~68 .sum_lutc_input = "datac";

dffeas \D_iw[20] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[20]~68_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cycloneive_lcell_comb \E_src1[16]~10 (
	.dataa(\D_iw[20]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[16]~10_combout ),
	.cout());
defparam \E_src1[16]~10 .lut_mask = 16'hAACC;
defparam \E_src1[16]~10 .sum_lutc_input = "datac";

dffeas \E_src1[16] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[16]~10_combout ),
	.asdata(\F_pc_plus_one[14]~28_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

dffeas \E_shift_rot_result[16] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[16]~11_combout ),
	.asdata(\E_src1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[16] .is_wysiwyg = "true";
defparam \E_shift_rot_result[16] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[15]~12 (
	.dataa(\E_shift_rot_result[16]~q ),
	.datab(\E_shift_rot_result[14]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[15]~12_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[15]~12 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[15]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[19]~69 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_19),
	.datad(out_data_buffer_19),
	.cin(gnd),
	.combout(\F_iw[19]~69_combout ),
	.cout());
defparam \F_iw[19]~69 .lut_mask = 16'hFFFE;
defparam \F_iw[19]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[19]~70 (
	.dataa(\F_iw[19]~69_combout ),
	.datab(out_payload_3),
	.datac(src_payload),
	.datad(\D_iw[1]~2_combout ),
	.cin(gnd),
	.combout(\F_iw[19]~70_combout ),
	.cout());
defparam \F_iw[19]~70 .lut_mask = 16'hFEFF;
defparam \F_iw[19]~70 .sum_lutc_input = "datac";

dffeas \D_iw[19] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[19]~70_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

cycloneive_lcell_comb \E_src1[15]~11 (
	.dataa(\D_iw[19]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[15]~11_combout ),
	.cout());
defparam \E_src1[15]~11 .lut_mask = 16'hAACC;
defparam \E_src1[15]~11 .sum_lutc_input = "datac";

dffeas \E_src1[15] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[15]~11_combout ),
	.asdata(\F_pc_plus_one[13]~26_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

dffeas \E_shift_rot_result[15] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[15]~12_combout ),
	.asdata(\E_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[15] .is_wysiwyg = "true";
defparam \E_shift_rot_result[15] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[14]~13 (
	.dataa(\E_shift_rot_result[15]~q ),
	.datab(\E_shift_rot_result[13]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[14]~13_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[14]~13 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[14]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~71 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_18),
	.datad(out_data_buffer_18),
	.cin(gnd),
	.combout(\F_iw[18]~71_combout ),
	.cout());
defparam \F_iw[18]~71 .lut_mask = 16'hFFFE;
defparam \F_iw[18]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~72 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[18]~71_combout ),
	.datac(out_payload_2),
	.datad(src_payload),
	.cin(gnd),
	.combout(\F_iw[18]~72_combout ),
	.cout());
defparam \F_iw[18]~72 .lut_mask = 16'hFFFE;
defparam \F_iw[18]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~73 (
	.dataa(\F_iw[18]~72_combout ),
	.datab(\hbreak_req~0_combout ),
	.datac(gnd),
	.datad(hbreak_enabled1),
	.cin(gnd),
	.combout(\F_iw[18]~73_combout ),
	.cout());
defparam \F_iw[18]~73 .lut_mask = 16'hEEFF;
defparam \F_iw[18]~73 .sum_lutc_input = "datac";

dffeas \D_iw[18] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[18]~73_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cycloneive_lcell_comb \E_src1[14]~12 (
	.dataa(\D_iw[18]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[14]~12_combout ),
	.cout());
defparam \E_src1[14]~12 .lut_mask = 16'hAACC;
defparam \E_src1[14]~12 .sum_lutc_input = "datac";

dffeas \E_src1[14] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[14]~12_combout ),
	.asdata(\F_pc_plus_one[12]~24_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

dffeas \E_shift_rot_result[14] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[14]~13_combout ),
	.asdata(\E_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[14] .is_wysiwyg = "true";
defparam \E_shift_rot_result[14] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[13]~14 (
	.dataa(\E_shift_rot_result[14]~q ),
	.datab(\E_shift_rot_result[12]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[13]~14_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[13]~14 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[13]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~74 (
	.dataa(out_valid),
	.datab(src1_valid),
	.datac(av_readdata_pre_17),
	.datad(out_data_buffer_17),
	.cin(gnd),
	.combout(\F_iw[17]~74_combout ),
	.cout());
defparam \F_iw[17]~74 .lut_mask = 16'hFFFE;
defparam \F_iw[17]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~75 (
	.dataa(\D_iw[1]~2_combout ),
	.datab(\F_iw[17]~74_combout ),
	.datac(out_payload_1),
	.datad(src_payload),
	.cin(gnd),
	.combout(\F_iw[17]~75_combout ),
	.cout());
defparam \F_iw[17]~75 .lut_mask = 16'hFFFE;
defparam \F_iw[17]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~79 (
	.dataa(\D_iw[1]~1_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\F_iw[17]~75_combout ),
	.cin(gnd),
	.combout(\F_iw[17]~79_combout ),
	.cout());
defparam \F_iw[17]~79 .lut_mask = 16'hFFDF;
defparam \F_iw[17]~79 .sum_lutc_input = "datac";

dffeas \D_iw[17] (
	.clk(wire_pll7_clk_0),
	.d(\F_iw[17]~79_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cycloneive_lcell_comb \E_src1[13]~13 (
	.dataa(\D_iw[17]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[13]~13_combout ),
	.cout());
defparam \E_src1[13]~13 .lut_mask = 16'hAACC;
defparam \E_src1[13]~13 .sum_lutc_input = "datac";

dffeas \E_src1[13] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[13]~13_combout ),
	.asdata(\F_pc_plus_one[11]~22_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

dffeas \E_shift_rot_result[13] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[13]~14_combout ),
	.asdata(\E_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[13] .is_wysiwyg = "true";
defparam \E_shift_rot_result[13] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[12]~15 (
	.dataa(\E_shift_rot_result[13]~q ),
	.datab(\E_shift_rot_result[11]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[12]~15_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[12]~15 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[12]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[12]~14 (
	.dataa(\D_iw[16]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[12]~14_combout ),
	.cout());
defparam \E_src1[12]~14 .lut_mask = 16'hAACC;
defparam \E_src1[12]~14 .sum_lutc_input = "datac";

dffeas \E_src1[12] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[12]~14_combout ),
	.asdata(\F_pc_plus_one[10]~20_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

dffeas \E_shift_rot_result[12] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[12]~15_combout ),
	.asdata(\E_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[12] .is_wysiwyg = "true";
defparam \E_shift_rot_result[12] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[11]~16 (
	.dataa(\E_shift_rot_result[12]~q ),
	.datab(\E_shift_rot_result[10]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[11]~16_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[11]~16 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[11]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[11]~15 (
	.dataa(\D_iw[15]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[11]~15_combout ),
	.cout());
defparam \E_src1[11]~15 .lut_mask = 16'hAACC;
defparam \E_src1[11]~15 .sum_lutc_input = "datac";

dffeas \E_src1[11] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[11]~15_combout ),
	.asdata(\F_pc_plus_one[9]~18_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

dffeas \E_shift_rot_result[11] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[11]~16_combout ),
	.asdata(\E_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[11] .is_wysiwyg = "true";
defparam \E_shift_rot_result[11] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[10]~17 (
	.dataa(\E_shift_rot_result[11]~q ),
	.datab(\E_shift_rot_result[9]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[10]~17_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[10]~17 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[10]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[10]~16 (
	.dataa(\D_iw[14]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[10]~16_combout ),
	.cout());
defparam \E_src1[10]~16 .lut_mask = 16'hAACC;
defparam \E_src1[10]~16 .sum_lutc_input = "datac";

dffeas \E_src1[10] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[10]~16_combout ),
	.asdata(\F_pc_plus_one[8]~16_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

dffeas \E_shift_rot_result[10] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[10]~17_combout ),
	.asdata(\E_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[10] .is_wysiwyg = "true";
defparam \E_shift_rot_result[10] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[9]~20 (
	.dataa(\E_shift_rot_result[10]~q ),
	.datab(\E_shift_rot_result[8]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[9]~20_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[9]~20 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[9]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[9]~17 (
	.dataa(\D_iw[13]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[9]~17_combout ),
	.cout());
defparam \E_src1[9]~17 .lut_mask = 16'hAACC;
defparam \E_src1[9]~17 .sum_lutc_input = "datac";

dffeas \E_src1[9] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[9]~17_combout ),
	.asdata(\F_pc_plus_one[7]~14_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

dffeas \E_shift_rot_result[9] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[9]~20_combout ),
	.asdata(\E_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[9] .is_wysiwyg = "true";
defparam \E_shift_rot_result[9] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[8]~21 (
	.dataa(\E_shift_rot_result[9]~q ),
	.datab(\E_shift_rot_result[7]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[8]~21_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[8]~21 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[8]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[8]~18 (
	.dataa(\D_iw[12]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[8]~18_combout ),
	.cout());
defparam \E_src1[8]~18 .lut_mask = 16'hAACC;
defparam \E_src1[8]~18 .sum_lutc_input = "datac";

dffeas \E_src1[8] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[8]~18_combout ),
	.asdata(\F_pc_plus_one[6]~12_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

dffeas \E_shift_rot_result[8] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[8]~21_combout ),
	.asdata(\E_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[8] .is_wysiwyg = "true";
defparam \E_shift_rot_result[8] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[7]~19 (
	.dataa(\E_shift_rot_result[8]~q ),
	.datab(\E_shift_rot_result[6]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[7]~19_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[7]~19 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[7]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[7]~19 (
	.dataa(\D_iw[11]~q ),
	.datab(\niosII_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(\R_src1~14_combout ),
	.cin(gnd),
	.combout(\E_src1[7]~19_combout ),
	.cout());
defparam \E_src1[7]~19 .lut_mask = 16'hAACC;
defparam \E_src1[7]~19 .sum_lutc_input = "datac";

dffeas \E_src1[7] (
	.clk(wire_pll7_clk_0),
	.d(\E_src1[7]~19_combout ),
	.asdata(\F_pc_plus_one[5]~10_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~15_combout ),
	.ena(vcc),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

dffeas \E_shift_rot_result[7] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[7]~19_combout ),
	.asdata(\E_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[7] .is_wysiwyg = "true";
defparam \E_shift_rot_result[7] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[6]~0 (
	.dataa(\E_shift_rot_result[7]~q ),
	.datab(\E_shift_rot_result[5]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[6]~0_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[6]~0 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[6]~0 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[6] (
	.clk(wire_pll7_clk_0),
	.d(\E_shift_rot_result_nxt[6]~0_combout ),
	.asdata(\E_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[6] .is_wysiwyg = "true";
defparam \E_shift_rot_result[6] .power_up = "low";

cycloneive_lcell_comb D_op_rdctl(
	.dataa(\Equal0~8_combout ),
	.datab(\Equal62~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_rdctl~combout ),
	.cout());
defparam D_op_rdctl.lut_mask = 16'hEFFF;
defparam D_op_rdctl.sum_lutc_input = "datac";

dffeas R_ctrl_rd_ctl_reg(
	.clk(wire_pll7_clk_0),
	.d(\D_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rd_ctl_reg~q ),
	.prn(vcc));
defparam R_ctrl_rd_ctl_reg.is_wysiwyg = "true";
defparam R_ctrl_rd_ctl_reg.power_up = "low";

cycloneive_lcell_comb \Equal0~6 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
defparam \Equal0~6 .lut_mask = 16'hF7FF;
defparam \Equal0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~2 (
	.dataa(\Equal0~6_combout ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~3_combout ),
	.datad(\D_ctrl_jmp_direct~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~2_combout ),
	.cout());
defparam \D_ctrl_br_cmp~2 .lut_mask = 16'hEFFF;
defparam \D_ctrl_br_cmp~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~5 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~5_combout ),
	.cout());
defparam \D_ctrl_br_cmp~5 .lut_mask = 16'hF7B3;
defparam \D_ctrl_br_cmp~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~3 (
	.dataa(\R_ctrl_br_nxt~1_combout ),
	.datab(\Equal0~8_combout ),
	.datac(\D_ctrl_br_cmp~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~3_combout ),
	.cout());
defparam \D_ctrl_br_cmp~3 .lut_mask = 16'hFEFE;
defparam \D_ctrl_br_cmp~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~4 (
	.dataa(\D_ctrl_br_cmp~2_combout ),
	.datab(\D_ctrl_br_cmp~3_combout ),
	.datac(\Equal62~0_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~4_combout ),
	.cout());
defparam \D_ctrl_br_cmp~4 .lut_mask = 16'hFFFE;
defparam \D_ctrl_br_cmp~4 .sum_lutc_input = "datac";

dffeas R_ctrl_br_cmp(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_br_cmp~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_cmp~q ),
	.prn(vcc));
defparam R_ctrl_br_cmp.is_wysiwyg = "true";
defparam R_ctrl_br_cmp.power_up = "low";

cycloneive_lcell_comb \E_alu_result~0 (
	.dataa(\R_ctrl_rd_ctl_reg~q ),
	.datab(\R_ctrl_br_cmp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_alu_result~0_combout ),
	.cout());
defparam \E_alu_result~0 .lut_mask = 16'hEEEE;
defparam \E_alu_result~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[26]~0 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[26]~0_combout ),
	.cout());
defparam \E_src2[26]~0 .lut_mask = 16'hAACC;
defparam \E_src2[26]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~2 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~6_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~2 .lut_mask = 16'hFAFC;
defparam \D_ctrl_unsigned_lo_imm16~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~3 (
	.dataa(\D_ctrl_unsigned_lo_imm16~1_combout ),
	.datab(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~3 .lut_mask = 16'hEFFF;
defparam \D_ctrl_unsigned_lo_imm16~3 .sum_lutc_input = "datac";

dffeas R_ctrl_unsigned_lo_imm16(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam R_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam R_ctrl_unsigned_lo_imm16.power_up = "low";

cycloneive_lcell_comb \R_src2_hi~0 (
	.dataa(\R_ctrl_force_src2_zero~q ),
	.datab(\R_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\R_src2_hi~0_combout ),
	.cout());
defparam \R_src2_hi~0 .lut_mask = 16'hEEEE;
defparam \R_src2_hi~0 .sum_lutc_input = "datac";

dffeas \E_src2[26] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[26]~0_combout ),
	.asdata(\D_iw[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cycloneive_lcell_comb \Add1~23 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[26]~q ),
	.cin(gnd),
	.combout(\Add1~23_combout ),
	.cout());
defparam \Add1~23 .lut_mask = 16'h0FF0;
defparam \Add1~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[25]~1 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[25]~1_combout ),
	.cout());
defparam \E_src2[25]~1 .lut_mask = 16'hAACC;
defparam \E_src2[25]~1 .sum_lutc_input = "datac";

dffeas \E_src2[25] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[25]~1_combout ),
	.asdata(\D_iw[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cycloneive_lcell_comb \Add1~24 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[25]~q ),
	.cin(gnd),
	.combout(\Add1~24_combout ),
	.cout());
defparam \Add1~24 .lut_mask = 16'h0FF0;
defparam \Add1~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[24]~2 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[24]~2_combout ),
	.cout());
defparam \E_src2[24]~2 .lut_mask = 16'hAACC;
defparam \E_src2[24]~2 .sum_lutc_input = "datac";

dffeas \E_src2[24] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[24]~2_combout ),
	.asdata(\D_iw[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cycloneive_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[24]~q ),
	.cin(gnd),
	.combout(\Add1~25_combout ),
	.cout());
defparam \Add1~25 .lut_mask = 16'h0FF0;
defparam \Add1~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[23]~3 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[23]~3_combout ),
	.cout());
defparam \E_src2[23]~3 .lut_mask = 16'hAACC;
defparam \E_src2[23]~3 .sum_lutc_input = "datac";

dffeas \E_src2[23] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[23]~3_combout ),
	.asdata(\D_iw[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cycloneive_lcell_comb \Add1~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[23]~q ),
	.cin(gnd),
	.combout(\Add1~26_combout ),
	.cout());
defparam \Add1~26 .lut_mask = 16'h0FF0;
defparam \Add1~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[22]~4 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[22]~4_combout ),
	.cout());
defparam \E_src2[22]~4 .lut_mask = 16'hAACC;
defparam \E_src2[22]~4 .sum_lutc_input = "datac";

dffeas \E_src2[22] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[22]~4_combout ),
	.asdata(\D_iw[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cycloneive_lcell_comb \Add1~27 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[22]~q ),
	.cin(gnd),
	.combout(\Add1~27_combout ),
	.cout());
defparam \Add1~27 .lut_mask = 16'h0FF0;
defparam \Add1~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[21]~5 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[21]~5_combout ),
	.cout());
defparam \E_src2[21]~5 .lut_mask = 16'hAACC;
defparam \E_src2[21]~5 .sum_lutc_input = "datac";

dffeas \E_src2[21] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[21]~5_combout ),
	.asdata(\D_iw[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cycloneive_lcell_comb \Add1~28 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[21]~q ),
	.cin(gnd),
	.combout(\Add1~28_combout ),
	.cout());
defparam \Add1~28 .lut_mask = 16'h0FF0;
defparam \Add1~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[20]~6 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[20]~6_combout ),
	.cout());
defparam \E_src2[20]~6 .lut_mask = 16'hAACC;
defparam \E_src2[20]~6 .sum_lutc_input = "datac";

dffeas \E_src2[20] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[20]~6_combout ),
	.asdata(\D_iw[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cycloneive_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[20]~q ),
	.cin(gnd),
	.combout(\Add1~29_combout ),
	.cout());
defparam \Add1~29 .lut_mask = 16'h0FF0;
defparam \Add1~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[19]~7 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[19]~7_combout ),
	.cout());
defparam \E_src2[19]~7 .lut_mask = 16'hAACC;
defparam \E_src2[19]~7 .sum_lutc_input = "datac";

dffeas \E_src2[19] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[19]~7_combout ),
	.asdata(\D_iw[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cycloneive_lcell_comb \Add1~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[19]~q ),
	.cin(gnd),
	.combout(\Add1~30_combout ),
	.cout());
defparam \Add1~30 .lut_mask = 16'h0FF0;
defparam \Add1~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[18]~8 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[18]~8_combout ),
	.cout());
defparam \E_src2[18]~8 .lut_mask = 16'hAACC;
defparam \E_src2[18]~8 .sum_lutc_input = "datac";

dffeas \E_src2[18] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[18]~8_combout ),
	.asdata(\D_iw[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cycloneive_lcell_comb \Add1~31 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[18]~q ),
	.cin(gnd),
	.combout(\Add1~31_combout ),
	.cout());
defparam \Add1~31 .lut_mask = 16'h0FF0;
defparam \Add1~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[17]~9 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[17]~9_combout ),
	.cout());
defparam \E_src2[17]~9 .lut_mask = 16'hAACC;
defparam \E_src2[17]~9 .sum_lutc_input = "datac";

dffeas \E_src2[17] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[17]~9_combout ),
	.asdata(\D_iw[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cycloneive_lcell_comb \Add1~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[17]~q ),
	.cin(gnd),
	.combout(\Add1~32_combout ),
	.cout());
defparam \Add1~32 .lut_mask = 16'h0FF0;
defparam \Add1~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[16]~10 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[16]~10_combout ),
	.cout());
defparam \E_src2[16]~10 .lut_mask = 16'hAACC;
defparam \E_src2[16]~10 .sum_lutc_input = "datac";

dffeas \E_src2[16] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[16]~10_combout ),
	.asdata(\D_iw[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

cycloneive_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[16]~q ),
	.cin(gnd),
	.combout(\Add1~33_combout ),
	.cout());
defparam \Add1~33 .lut_mask = 16'h0FF0;
defparam \Add1~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[15]~9 (
	.dataa(\D_iw[21]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[15]~9_combout ),
	.cout());
defparam \R_src2_lo[15]~9 .lut_mask = 16'hACFF;
defparam \R_src2_lo[15]~9 .sum_lutc_input = "datac";

dffeas \E_src2[15] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[15]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

cycloneive_lcell_comb \Add1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[15]~q ),
	.cin(gnd),
	.combout(\Add1~34_combout ),
	.cout());
defparam \Add1~34 .lut_mask = 16'h0FF0;
defparam \Add1~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[14]~10 (
	.dataa(\D_iw[20]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[14]~10_combout ),
	.cout());
defparam \R_src2_lo[14]~10 .lut_mask = 16'hACFF;
defparam \R_src2_lo[14]~10 .sum_lutc_input = "datac";

dffeas \E_src2[14] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[14]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

cycloneive_lcell_comb \Add1~35 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[14]~q ),
	.cin(gnd),
	.combout(\Add1~35_combout ),
	.cout());
defparam \Add1~35 .lut_mask = 16'h0FF0;
defparam \Add1~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[13]~11 (
	.dataa(\D_iw[19]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[13]~11_combout ),
	.cout());
defparam \R_src2_lo[13]~11 .lut_mask = 16'hACFF;
defparam \R_src2_lo[13]~11 .sum_lutc_input = "datac";

dffeas \E_src2[13] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[13]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

cycloneive_lcell_comb \Add1~36 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[13]~q ),
	.cin(gnd),
	.combout(\Add1~36_combout ),
	.cout());
defparam \Add1~36 .lut_mask = 16'h0FF0;
defparam \Add1~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[12]~12 (
	.dataa(\D_iw[18]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[12]~12_combout ),
	.cout());
defparam \R_src2_lo[12]~12 .lut_mask = 16'hACFF;
defparam \R_src2_lo[12]~12 .sum_lutc_input = "datac";

dffeas \E_src2[12] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[12]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

cycloneive_lcell_comb \Add1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[12]~q ),
	.cin(gnd),
	.combout(\Add1~37_combout ),
	.cout());
defparam \Add1~37 .lut_mask = 16'h0FF0;
defparam \Add1~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[11]~13 (
	.dataa(\D_iw[17]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[11]~13_combout ),
	.cout());
defparam \R_src2_lo[11]~13 .lut_mask = 16'hACFF;
defparam \R_src2_lo[11]~13 .sum_lutc_input = "datac";

dffeas \E_src2[11] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[11]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

cycloneive_lcell_comb \Add1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[11]~q ),
	.cin(gnd),
	.combout(\Add1~38_combout ),
	.cout());
defparam \Add1~38 .lut_mask = 16'h0FF0;
defparam \Add1~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[10]~14 (
	.dataa(\D_iw[16]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[10]~14_combout ),
	.cout());
defparam \R_src2_lo[10]~14 .lut_mask = 16'hACFF;
defparam \R_src2_lo[10]~14 .sum_lutc_input = "datac";

dffeas \E_src2[10] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[10]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

cycloneive_lcell_comb \Add1~39 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[10]~q ),
	.cin(gnd),
	.combout(\Add1~39_combout ),
	.cout());
defparam \Add1~39 .lut_mask = 16'h0FF0;
defparam \Add1~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[9]~15 (
	.dataa(\D_iw[15]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[9]~15_combout ),
	.cout());
defparam \R_src2_lo[9]~15 .lut_mask = 16'hACFF;
defparam \R_src2_lo[9]~15 .sum_lutc_input = "datac";

dffeas \E_src2[9] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[9]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

cycloneive_lcell_comb \Add1~40 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[9]~q ),
	.cin(gnd),
	.combout(\Add1~40_combout ),
	.cout());
defparam \Add1~40 .lut_mask = 16'h0FF0;
defparam \Add1~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[8]~16 (
	.dataa(\D_iw[14]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[8]~16_combout ),
	.cout());
defparam \R_src2_lo[8]~16 .lut_mask = 16'hACFF;
defparam \R_src2_lo[8]~16 .sum_lutc_input = "datac";

dffeas \E_src2[8] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[8]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

cycloneive_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[8]~q ),
	.cin(gnd),
	.combout(\Add1~41_combout ),
	.cout());
defparam \Add1~41 .lut_mask = 16'h0FF0;
defparam \Add1~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[7]~17 (
	.dataa(\D_iw[13]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[7]~17_combout ),
	.cout());
defparam \R_src2_lo[7]~17 .lut_mask = 16'hACFF;
defparam \R_src2_lo[7]~17 .sum_lutc_input = "datac";

dffeas \E_src2[7] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_lo[7]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

cycloneive_lcell_comb \Add1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[7]~q ),
	.cin(gnd),
	.combout(\Add1~42_combout ),
	.cout());
defparam \Add1~42 .lut_mask = 16'h0FF0;
defparam \Add1~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~43 (
	.dataa(\Add1~42_combout ),
	.datab(\E_src1[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~22 ),
	.combout(\Add1~43_combout ),
	.cout(\Add1~44 ));
defparam \Add1~43 .lut_mask = 16'h96EF;
defparam \Add1~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~45 (
	.dataa(\Add1~41_combout ),
	.datab(\E_src1[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~44 ),
	.combout(\Add1~45_combout ),
	.cout(\Add1~46 ));
defparam \Add1~45 .lut_mask = 16'h967F;
defparam \Add1~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~47 (
	.dataa(\Add1~40_combout ),
	.datab(\E_src1[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~46 ),
	.combout(\Add1~47_combout ),
	.cout(\Add1~48 ));
defparam \Add1~47 .lut_mask = 16'h96EF;
defparam \Add1~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~49 (
	.dataa(\Add1~39_combout ),
	.datab(\E_src1[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~48 ),
	.combout(\Add1~49_combout ),
	.cout(\Add1~50 ));
defparam \Add1~49 .lut_mask = 16'h967F;
defparam \Add1~49 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~51 (
	.dataa(\Add1~38_combout ),
	.datab(\E_src1[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~50 ),
	.combout(\Add1~51_combout ),
	.cout(\Add1~52 ));
defparam \Add1~51 .lut_mask = 16'h96EF;
defparam \Add1~51 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~53 (
	.dataa(\Add1~37_combout ),
	.datab(\E_src1[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~52 ),
	.combout(\Add1~53_combout ),
	.cout(\Add1~54 ));
defparam \Add1~53 .lut_mask = 16'h967F;
defparam \Add1~53 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~55 (
	.dataa(\Add1~36_combout ),
	.datab(\E_src1[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~54 ),
	.combout(\Add1~55_combout ),
	.cout(\Add1~56 ));
defparam \Add1~55 .lut_mask = 16'h96EF;
defparam \Add1~55 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~57 (
	.dataa(\Add1~35_combout ),
	.datab(\E_src1[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~56 ),
	.combout(\Add1~57_combout ),
	.cout(\Add1~58 ));
defparam \Add1~57 .lut_mask = 16'h967F;
defparam \Add1~57 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~59 (
	.dataa(\Add1~34_combout ),
	.datab(\E_src1[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~58 ),
	.combout(\Add1~59_combout ),
	.cout(\Add1~60 ));
defparam \Add1~59 .lut_mask = 16'h96EF;
defparam \Add1~59 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~61 (
	.dataa(\Add1~33_combout ),
	.datab(\E_src1[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~60 ),
	.combout(\Add1~61_combout ),
	.cout(\Add1~62 ));
defparam \Add1~61 .lut_mask = 16'h967F;
defparam \Add1~61 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~63 (
	.dataa(\Add1~32_combout ),
	.datab(\E_src1[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~62 ),
	.combout(\Add1~63_combout ),
	.cout(\Add1~64 ));
defparam \Add1~63 .lut_mask = 16'h96EF;
defparam \Add1~63 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~65 (
	.dataa(\Add1~31_combout ),
	.datab(\E_src1[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~64 ),
	.combout(\Add1~65_combout ),
	.cout(\Add1~66 ));
defparam \Add1~65 .lut_mask = 16'h967F;
defparam \Add1~65 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~67 (
	.dataa(\Add1~30_combout ),
	.datab(\E_src1[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~66 ),
	.combout(\Add1~67_combout ),
	.cout(\Add1~68 ));
defparam \Add1~67 .lut_mask = 16'h96EF;
defparam \Add1~67 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~69 (
	.dataa(\Add1~29_combout ),
	.datab(\E_src1[20]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~68 ),
	.combout(\Add1~69_combout ),
	.cout(\Add1~70 ));
defparam \Add1~69 .lut_mask = 16'h967F;
defparam \Add1~69 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~71 (
	.dataa(\Add1~28_combout ),
	.datab(\E_src1[21]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~70 ),
	.combout(\Add1~71_combout ),
	.cout(\Add1~72 ));
defparam \Add1~71 .lut_mask = 16'h96EF;
defparam \Add1~71 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~73 (
	.dataa(\Add1~27_combout ),
	.datab(\E_src1[22]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~72 ),
	.combout(\Add1~73_combout ),
	.cout(\Add1~74 ));
defparam \Add1~73 .lut_mask = 16'h967F;
defparam \Add1~73 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~75 (
	.dataa(\Add1~26_combout ),
	.datab(\E_src1[23]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~74 ),
	.combout(\Add1~75_combout ),
	.cout(\Add1~76 ));
defparam \Add1~75 .lut_mask = 16'h96EF;
defparam \Add1~75 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~77 (
	.dataa(\Add1~25_combout ),
	.datab(\E_src1[24]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~76 ),
	.combout(\Add1~77_combout ),
	.cout(\Add1~78 ));
defparam \Add1~77 .lut_mask = 16'h967F;
defparam \Add1~77 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~79 (
	.dataa(\Add1~24_combout ),
	.datab(\E_src1[25]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~78 ),
	.combout(\Add1~79_combout ),
	.cout(\Add1~80 ));
defparam \Add1~79 .lut_mask = 16'h96EF;
defparam \Add1~79 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~81 (
	.dataa(\Add1~23_combout ),
	.datab(\E_src1[26]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~80 ),
	.combout(\Add1~81_combout ),
	.cout(\Add1~82 ));
defparam \Add1~81 .lut_mask = 16'h967F;
defparam \Add1~81 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_logic_result[26]~1 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[26]~q ),
	.datac(\E_src1[26]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[26]~1_combout ),
	.cout());
defparam \E_logic_result[26]~1 .lut_mask = 16'h6996;
defparam \E_logic_result[26]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[26]~0 (
	.dataa(\Add1~81_combout ),
	.datab(\E_logic_result[26]~1_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[26]~0_combout ),
	.cout());
defparam \W_alu_result[26]~0 .lut_mask = 16'hAACC;
defparam \W_alu_result[26]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[25]~2 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[25]~q ),
	.datac(\E_src1[25]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[25]~2_combout ),
	.cout());
defparam \E_logic_result[25]~2 .lut_mask = 16'h6996;
defparam \E_logic_result[25]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[25]~1 (
	.dataa(\Add1~79_combout ),
	.datab(\E_logic_result[25]~2_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[25]~1_combout ),
	.cout());
defparam \W_alu_result[25]~1 .lut_mask = 16'hAACC;
defparam \W_alu_result[25]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[24]~3 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[24]~q ),
	.datac(\E_src1[24]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[24]~3_combout ),
	.cout());
defparam \E_logic_result[24]~3 .lut_mask = 16'h6996;
defparam \E_logic_result[24]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[24]~2 (
	.dataa(\Add1~77_combout ),
	.datab(\E_logic_result[24]~3_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[24]~2_combout ),
	.cout());
defparam \W_alu_result[24]~2 .lut_mask = 16'hAACC;
defparam \W_alu_result[24]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[23]~4 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[23]~q ),
	.datac(\E_src1[23]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[23]~4_combout ),
	.cout());
defparam \E_logic_result[23]~4 .lut_mask = 16'h6996;
defparam \E_logic_result[23]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[23]~3 (
	.dataa(\Add1~75_combout ),
	.datab(\E_logic_result[23]~4_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[23]~3_combout ),
	.cout());
defparam \W_alu_result[23]~3 .lut_mask = 16'hAACC;
defparam \W_alu_result[23]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[22]~5 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[22]~q ),
	.datac(\E_src1[22]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[22]~5_combout ),
	.cout());
defparam \E_logic_result[22]~5 .lut_mask = 16'h6996;
defparam \E_logic_result[22]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[22]~4 (
	.dataa(\Add1~73_combout ),
	.datab(\E_logic_result[22]~5_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[22]~4_combout ),
	.cout());
defparam \W_alu_result[22]~4 .lut_mask = 16'hAACC;
defparam \W_alu_result[22]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[21]~6 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[21]~q ),
	.datac(\E_src1[21]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[21]~6_combout ),
	.cout());
defparam \E_logic_result[21]~6 .lut_mask = 16'h6996;
defparam \E_logic_result[21]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[21]~5 (
	.dataa(\Add1~71_combout ),
	.datab(\E_logic_result[21]~6_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[21]~5_combout ),
	.cout());
defparam \W_alu_result[21]~5 .lut_mask = 16'hAACC;
defparam \W_alu_result[21]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[20]~7 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[20]~q ),
	.datac(\E_src1[20]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[20]~7_combout ),
	.cout());
defparam \E_logic_result[20]~7 .lut_mask = 16'h6996;
defparam \E_logic_result[20]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[20]~6 (
	.dataa(\Add1~69_combout ),
	.datab(\E_logic_result[20]~7_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[20]~6_combout ),
	.cout());
defparam \W_alu_result[20]~6 .lut_mask = 16'hAACC;
defparam \W_alu_result[20]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[19]~8 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[19]~q ),
	.datac(\E_src1[19]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[19]~8_combout ),
	.cout());
defparam \E_logic_result[19]~8 .lut_mask = 16'h6996;
defparam \E_logic_result[19]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[19]~7 (
	.dataa(\Add1~67_combout ),
	.datab(\E_logic_result[19]~8_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[19]~7_combout ),
	.cout());
defparam \W_alu_result[19]~7 .lut_mask = 16'hAACC;
defparam \W_alu_result[19]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[18]~9 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[18]~q ),
	.datac(\E_src1[18]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[18]~9_combout ),
	.cout());
defparam \E_logic_result[18]~9 .lut_mask = 16'h6996;
defparam \E_logic_result[18]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[18]~8 (
	.dataa(\Add1~65_combout ),
	.datab(\E_logic_result[18]~9_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[18]~8_combout ),
	.cout());
defparam \W_alu_result[18]~8 .lut_mask = 16'hAACC;
defparam \W_alu_result[18]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[17]~10 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[17]~q ),
	.datac(\E_src1[17]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[17]~10_combout ),
	.cout());
defparam \E_logic_result[17]~10 .lut_mask = 16'h6996;
defparam \E_logic_result[17]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[17]~9 (
	.dataa(\Add1~63_combout ),
	.datab(\E_logic_result[17]~10_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[17]~9_combout ),
	.cout());
defparam \W_alu_result[17]~9 .lut_mask = 16'hAACC;
defparam \W_alu_result[17]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[16]~11 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[16]~q ),
	.datac(\E_src1[16]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[16]~11_combout ),
	.cout());
defparam \E_logic_result[16]~11 .lut_mask = 16'h6996;
defparam \E_logic_result[16]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[16]~10 (
	.dataa(\Add1~61_combout ),
	.datab(\E_logic_result[16]~11_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[16]~10_combout ),
	.cout());
defparam \W_alu_result[16]~10 .lut_mask = 16'hAACC;
defparam \W_alu_result[16]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[15]~12 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[15]~q ),
	.datac(\E_src1[15]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[15]~12_combout ),
	.cout());
defparam \E_logic_result[15]~12 .lut_mask = 16'h6996;
defparam \E_logic_result[15]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[15]~11 (
	.dataa(\Add1~59_combout ),
	.datab(\E_logic_result[15]~12_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[15]~11_combout ),
	.cout());
defparam \W_alu_result[15]~11 .lut_mask = 16'hAACC;
defparam \W_alu_result[15]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[14]~13 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[14]~q ),
	.datac(\E_src1[14]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[14]~13_combout ),
	.cout());
defparam \E_logic_result[14]~13 .lut_mask = 16'h6996;
defparam \E_logic_result[14]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[14]~12 (
	.dataa(\Add1~57_combout ),
	.datab(\E_logic_result[14]~13_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[14]~12_combout ),
	.cout());
defparam \W_alu_result[14]~12 .lut_mask = 16'hAACC;
defparam \W_alu_result[14]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[13]~14 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[13]~q ),
	.datac(\E_src1[13]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[13]~14_combout ),
	.cout());
defparam \E_logic_result[13]~14 .lut_mask = 16'h6996;
defparam \E_logic_result[13]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[13]~13 (
	.dataa(\Add1~55_combout ),
	.datab(\E_logic_result[13]~14_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[13]~13_combout ),
	.cout());
defparam \W_alu_result[13]~13 .lut_mask = 16'hAACC;
defparam \W_alu_result[13]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[12]~15 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[12]~q ),
	.datac(\E_src1[12]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[12]~15_combout ),
	.cout());
defparam \E_logic_result[12]~15 .lut_mask = 16'h6996;
defparam \E_logic_result[12]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[12]~14 (
	.dataa(\Add1~53_combout ),
	.datab(\E_logic_result[12]~15_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[12]~14_combout ),
	.cout());
defparam \W_alu_result[12]~14 .lut_mask = 16'hAACC;
defparam \W_alu_result[12]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[11]~16 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[11]~q ),
	.datac(\E_src1[11]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[11]~16_combout ),
	.cout());
defparam \E_logic_result[11]~16 .lut_mask = 16'h6996;
defparam \E_logic_result[11]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[11]~15 (
	.dataa(\Add1~51_combout ),
	.datab(\E_logic_result[11]~16_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[11]~15_combout ),
	.cout());
defparam \W_alu_result[11]~15 .lut_mask = 16'hAACC;
defparam \W_alu_result[11]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[10]~17 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[10]~q ),
	.datac(\E_src1[10]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[10]~17_combout ),
	.cout());
defparam \E_logic_result[10]~17 .lut_mask = 16'h6996;
defparam \E_logic_result[10]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[10]~16 (
	.dataa(\Add1~49_combout ),
	.datab(\E_logic_result[10]~17_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[10]~16_combout ),
	.cout());
defparam \W_alu_result[10]~16 .lut_mask = 16'hAACC;
defparam \W_alu_result[10]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[5]~18 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[5]~q ),
	.datac(\E_src1[5]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[5]~18_combout ),
	.cout());
defparam \E_logic_result[5]~18 .lut_mask = 16'h6996;
defparam \E_logic_result[5]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[5]~21 (
	.dataa(\Add1~19_combout ),
	.datab(\E_logic_result[5]~18_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[5]~21_combout ),
	.cout());
defparam \W_alu_result[5]~21 .lut_mask = 16'hAACC;
defparam \W_alu_result[5]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[7]~19 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[7]~q ),
	.datac(\E_src1[7]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[7]~19_combout ),
	.cout());
defparam \E_logic_result[7]~19 .lut_mask = 16'h6996;
defparam \E_logic_result[7]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[7]~19 (
	.dataa(\Add1~43_combout ),
	.datab(\E_logic_result[7]~19_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[7]~19_combout ),
	.cout());
defparam \W_alu_result[7]~19 .lut_mask = 16'hAACC;
defparam \W_alu_result[7]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[9]~20 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[9]~q ),
	.datac(\E_src1[9]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[9]~20_combout ),
	.cout());
defparam \E_logic_result[9]~20 .lut_mask = 16'h6996;
defparam \E_logic_result[9]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[9]~17 (
	.dataa(\Add1~47_combout ),
	.datab(\E_logic_result[9]~20_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[9]~17_combout ),
	.cout());
defparam \W_alu_result[9]~17 .lut_mask = 16'hAACC;
defparam \W_alu_result[9]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[8]~21 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[8]~q ),
	.datac(\E_src1[8]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[8]~21_combout ),
	.cout());
defparam \E_logic_result[8]~21 .lut_mask = 16'h6996;
defparam \E_logic_result[8]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[8]~18 (
	.dataa(\Add1~45_combout ),
	.datab(\E_logic_result[8]~21_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[8]~18_combout ),
	.cout());
defparam \W_alu_result[8]~18 .lut_mask = 16'hAACC;
defparam \W_alu_result[8]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[4]~22 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[4]~q ),
	.datac(\E_src1[4]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[4]~22_combout ),
	.cout());
defparam \E_logic_result[4]~22 .lut_mask = 16'h6996;
defparam \E_logic_result[4]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[4]~22 (
	.dataa(\Add1~17_combout ),
	.datab(\E_logic_result[4]~22_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[4]~22_combout ),
	.cout());
defparam \W_alu_result[4]~22 .lut_mask = 16'hAACC;
defparam \W_alu_result[4]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[3]~23 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[3]~q ),
	.datac(\E_src1[3]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[3]~23_combout ),
	.cout());
defparam \E_logic_result[3]~23 .lut_mask = 16'h6996;
defparam \E_logic_result[3]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[3]~23 (
	.dataa(\Add1~15_combout ),
	.datab(\E_logic_result[3]~23_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[3]~23_combout ),
	.cout());
defparam \W_alu_result[3]~23 .lut_mask = 16'hAACC;
defparam \W_alu_result[3]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[2]~24 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[2]~q ),
	.datac(\E_src1[2]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[2]~24_combout ),
	.cout());
defparam \E_logic_result[2]~24 .lut_mask = 16'h6996;
defparam \E_logic_result[2]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[2]~24 (
	.dataa(\Add1~13_combout ),
	.datab(\E_logic_result[2]~24_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[2]~24_combout ),
	.cout());
defparam \W_alu_result[2]~24 .lut_mask = 16'hAACC;
defparam \W_alu_result[2]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[24]~0 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[24]~0_combout ),
	.cout());
defparam \d_writedata[24]~0 .lut_mask = 16'hAACC;
defparam \d_writedata[24]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem8~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~0_combout ),
	.cout());
defparam \D_ctrl_mem8~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem8~1 (
	.dataa(\D_ctrl_mem8~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~1_combout ),
	.cout());
defparam \D_ctrl_mem8~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[25]~1 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[25]~1_combout ),
	.cout());
defparam \d_writedata[25]~1 .lut_mask = 16'hAACC;
defparam \d_writedata[25]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[26]~2 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[26]~2_combout ),
	.cout());
defparam \d_writedata[26]~2 .lut_mask = 16'hAACC;
defparam \d_writedata[26]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[27]~3 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[27]~3_combout ),
	.cout());
defparam \d_writedata[27]~3 .lut_mask = 16'hAACC;
defparam \d_writedata[27]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[28]~4 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[28]~4_combout ),
	.cout());
defparam \d_writedata[28]~4 .lut_mask = 16'hAACC;
defparam \d_writedata[28]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[29]~5 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[29]~5_combout ),
	.cout());
defparam \d_writedata[29]~5 .lut_mask = 16'hAACC;
defparam \d_writedata[29]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[30]~6 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[30]~6_combout ),
	.cout());
defparam \d_writedata[30]~6 .lut_mask = 16'hAACC;
defparam \d_writedata[30]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[31]~7 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[31]~7_combout ),
	.cout());
defparam \d_writedata[31]~7 .lut_mask = 16'hAACC;
defparam \d_writedata[31]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb d_read_nxt(
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(d_read1),
	.datad(WideOr1),
	.cin(gnd),
	.combout(\d_read_nxt~combout ),
	.cout());
defparam d_read_nxt.lut_mask = 16'hFFFE;
defparam d_read_nxt.sum_lutc_input = "datac";

cycloneive_lcell_comb E_st_stall(
	.dataa(d_write1),
	.datab(\E_new_inst~q ),
	.datac(\R_ctrl_st~q ),
	.datad(av_waitrequest),
	.cin(gnd),
	.combout(\E_st_stall~combout ),
	.cout());
defparam E_st_stall.lut_mask = 16'hFFFE;
defparam E_st_stall.sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[0]~0 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~9_combout ),
	.datad(\Add1~11_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[0]~0_combout ),
	.cout());
defparam \E_mem_byte_en[0]~0 .lut_mask = 16'h6FFF;
defparam \E_mem_byte_en[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[1]~1 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~9_combout ),
	.datad(\Add1~11_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[1]~1_combout ),
	.cout());
defparam \E_mem_byte_en[1]~1 .lut_mask = 16'hF6FF;
defparam \E_mem_byte_en[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_read_nxt~0 (
	.dataa(\W_valid~q ),
	.datab(read_accepted),
	.datac(i_read1),
	.datad(src1_valid1),
	.cin(gnd),
	.combout(\i_read_nxt~0_combout ),
	.cout());
defparam \i_read_nxt~0 .lut_mask = 16'hFFF7;
defparam \i_read_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~0 (
	.dataa(\Equal0~8_combout ),
	.datab(\Equal62~8_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~0_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_uncond_cti_non_br~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~2 (
	.dataa(\D_ctrl_jmp_direct~1_combout ),
	.datab(\D_ctrl_uncond_cti_non_br~0_combout ),
	.datac(gnd),
	.datad(\D_ctrl_uncond_cti_non_br~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~2_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~2 .lut_mask = 16'hEEFF;
defparam \D_ctrl_uncond_cti_non_br~2 .sum_lutc_input = "datac";

dffeas R_ctrl_uncond_cti_non_br(
	.clk(wire_pll7_clk_0),
	.d(\D_ctrl_uncond_cti_non_br~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_uncond_cti_non_br~q ),
	.prn(vcc));
defparam R_ctrl_uncond_cti_non_br.is_wysiwyg = "true";
defparam R_ctrl_uncond_cti_non_br.power_up = "low";

cycloneive_lcell_comb \Equal0~20 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~20_combout ),
	.cout());
defparam \Equal0~20 .lut_mask = 16'hF7F7;
defparam \Equal0~20 .sum_lutc_input = "datac";

dffeas R_ctrl_br_uncond(
	.clk(wire_pll7_clk_0),
	.d(\Equal0~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_uncond~q ),
	.prn(vcc));
defparam R_ctrl_br_uncond.is_wysiwyg = "true";
defparam R_ctrl_br_uncond.power_up = "low";

dffeas \R_compare_op[1] (
	.clk(wire_pll7_clk_0),
	.d(\D_logic_op_raw[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[1]~q ),
	.prn(vcc));
defparam \R_compare_op[1] .is_wysiwyg = "true";
defparam \R_compare_op[1] .power_up = "low";

cycloneive_lcell_comb \D_logic_op_raw[0]~1 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\D_logic_op_raw[0]~1_combout ),
	.cout());
defparam \D_logic_op_raw[0]~1 .lut_mask = 16'hEFFE;
defparam \D_logic_op_raw[0]~1 .sum_lutc_input = "datac";

dffeas \R_compare_op[0] (
	.clk(wire_pll7_clk_0),
	.d(\D_logic_op_raw[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[0]~q ),
	.prn(vcc));
defparam \R_compare_op[0] .is_wysiwyg = "true";
defparam \R_compare_op[0] .power_up = "low";

cycloneive_lcell_comb \Equal127~0 (
	.dataa(\E_logic_result[26]~1_combout ),
	.datab(\E_logic_result[25]~2_combout ),
	.datac(\E_logic_result[24]~3_combout ),
	.datad(\E_logic_result[23]~4_combout ),
	.cin(gnd),
	.combout(\Equal127~0_combout ),
	.cout());
defparam \Equal127~0 .lut_mask = 16'h7FFF;
defparam \Equal127~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~1 (
	.dataa(\E_logic_result[22]~5_combout ),
	.datab(\E_logic_result[21]~6_combout ),
	.datac(\E_logic_result[20]~7_combout ),
	.datad(\E_logic_result[19]~8_combout ),
	.cin(gnd),
	.combout(\Equal127~1_combout ),
	.cout());
defparam \Equal127~1 .lut_mask = 16'h7FFF;
defparam \Equal127~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~2 (
	.dataa(\E_logic_result[18]~9_combout ),
	.datab(\E_logic_result[17]~10_combout ),
	.datac(\E_logic_result[16]~11_combout ),
	.datad(\E_logic_result[15]~12_combout ),
	.cin(gnd),
	.combout(\Equal127~2_combout ),
	.cout());
defparam \Equal127~2 .lut_mask = 16'h7FFF;
defparam \Equal127~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~3 (
	.dataa(\E_logic_result[14]~13_combout ),
	.datab(\E_logic_result[13]~14_combout ),
	.datac(\E_logic_result[12]~15_combout ),
	.datad(\E_logic_result[11]~16_combout ),
	.cin(gnd),
	.combout(\Equal127~3_combout ),
	.cout());
defparam \Equal127~3 .lut_mask = 16'h7FFF;
defparam \Equal127~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~4 (
	.dataa(\Equal127~0_combout ),
	.datab(\Equal127~1_combout ),
	.datac(\Equal127~2_combout ),
	.datad(\Equal127~3_combout ),
	.cin(gnd),
	.combout(\Equal127~4_combout ),
	.cout());
defparam \Equal127~4 .lut_mask = 16'hFFFE;
defparam \Equal127~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~5 (
	.dataa(\E_logic_result[7]~19_combout ),
	.datab(\E_logic_result[10]~17_combout ),
	.datac(\E_logic_result[9]~20_combout ),
	.datad(\E_logic_result[8]~21_combout ),
	.cin(gnd),
	.combout(\Equal127~5_combout ),
	.cout());
defparam \Equal127~5 .lut_mask = 16'h7FFF;
defparam \Equal127~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~6 (
	.dataa(\E_logic_result[5]~18_combout ),
	.datab(\E_logic_result[6]~0_combout ),
	.datac(\E_logic_result[4]~22_combout ),
	.datad(\E_logic_result[3]~23_combout ),
	.cin(gnd),
	.combout(\Equal127~6_combout ),
	.cout());
defparam \Equal127~6 .lut_mask = 16'h7FFF;
defparam \Equal127~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_hi[15]~1 (
	.dataa(\D_iw[21]~q ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datac(\R_ctrl_hi_imm16~q ),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~1_combout ),
	.cout());
defparam \R_src2_hi[15]~1 .lut_mask = 16'hEFFE;
defparam \R_src2_hi[15]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_hi[15]~2 (
	.dataa(\R_src2_hi[15]~1_combout ),
	.datab(gnd),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(\R_ctrl_unsigned_lo_imm16~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~2_combout ),
	.cout());
defparam \R_src2_hi[15]~2 .lut_mask = 16'hAFFF;
defparam \R_src2_hi[15]~2 .sum_lutc_input = "datac";

dffeas \E_src2[31] (
	.clk(wire_pll7_clk_0),
	.d(\R_src2_hi[15]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[31]~25 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_src1[31]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[31]~25_combout ),
	.cout());
defparam \E_logic_result[31]~25 .lut_mask = 16'h6996;
defparam \E_logic_result[31]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[30]~11 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[30]~11_combout ),
	.cout());
defparam \E_src2[30]~11 .lut_mask = 16'hAACC;
defparam \E_src2[30]~11 .sum_lutc_input = "datac";

dffeas \E_src2[30] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[30]~11_combout ),
	.asdata(\D_iw[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[30]~26 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[30]~q ),
	.datac(\E_src1[30]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[30]~26_combout ),
	.cout());
defparam \E_logic_result[30]~26 .lut_mask = 16'h6996;
defparam \E_logic_result[30]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[29]~12 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[29]~12_combout ),
	.cout());
defparam \E_src2[29]~12 .lut_mask = 16'hAACC;
defparam \E_src2[29]~12 .sum_lutc_input = "datac";

dffeas \E_src2[29] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[29]~12_combout ),
	.asdata(\D_iw[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[29]~27 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[29]~q ),
	.datac(\E_src1[29]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[29]~27_combout ),
	.cout());
defparam \E_logic_result[29]~27 .lut_mask = 16'h6996;
defparam \E_logic_result[29]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~7 (
	.dataa(\E_logic_result[2]~24_combout ),
	.datab(\E_logic_result[31]~25_combout ),
	.datac(\E_logic_result[30]~26_combout ),
	.datad(\E_logic_result[29]~27_combout ),
	.cin(gnd),
	.combout(\Equal127~7_combout ),
	.cout());
defparam \Equal127~7 .lut_mask = 16'h7FFF;
defparam \Equal127~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[28]~13 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[28]~13_combout ),
	.cout());
defparam \E_src2[28]~13 .lut_mask = 16'hAACC;
defparam \E_src2[28]~13 .sum_lutc_input = "datac";

dffeas \E_src2[28] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[28]~13_combout ),
	.asdata(\D_iw[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[28]~28 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[28]~q ),
	.datac(\E_src1[28]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[28]~28_combout ),
	.cout());
defparam \E_logic_result[28]~28 .lut_mask = 16'h6996;
defparam \E_logic_result[28]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[27]~14 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[27]~14_combout ),
	.cout());
defparam \E_src2[27]~14 .lut_mask = 16'hAACC;
defparam \E_src2[27]~14 .sum_lutc_input = "datac";

dffeas \E_src2[27] (
	.clk(wire_pll7_clk_0),
	.d(\E_src2[27]~14_combout ),
	.asdata(\D_iw[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[27]~29 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[27]~q ),
	.datac(\E_src1[27]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[27]~29_combout ),
	.cout());
defparam \E_logic_result[27]~29 .lut_mask = 16'h6996;
defparam \E_logic_result[27]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[1]~30 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[1]~q ),
	.datac(\E_src1[1]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[1]~30_combout ),
	.cout());
defparam \E_logic_result[1]~30 .lut_mask = 16'h6996;
defparam \E_logic_result[1]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[0]~31 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[0]~q ),
	.datac(\E_src1[0]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[0]~31_combout ),
	.cout());
defparam \E_logic_result[0]~31 .lut_mask = 16'h6996;
defparam \E_logic_result[0]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~8 (
	.dataa(\E_logic_result[28]~28_combout ),
	.datab(\E_logic_result[27]~29_combout ),
	.datac(\E_logic_result[1]~30_combout ),
	.datad(\E_logic_result[0]~31_combout ),
	.cin(gnd),
	.combout(\Equal127~8_combout ),
	.cout());
defparam \Equal127~8 .lut_mask = 16'h7FFF;
defparam \Equal127~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~9 (
	.dataa(\Equal127~5_combout ),
	.datab(\Equal127~6_combout ),
	.datac(\Equal127~7_combout ),
	.datad(\Equal127~8_combout ),
	.cin(gnd),
	.combout(\Equal127~9_combout ),
	.cout());
defparam \Equal127~9 .lut_mask = 16'hFFFE;
defparam \Equal127~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_cmp_result~0 (
	.dataa(\R_compare_op[1]~q ),
	.datab(\R_compare_op[0]~q ),
	.datac(\Equal127~4_combout ),
	.datad(\Equal127~9_combout ),
	.cin(gnd),
	.combout(\E_cmp_result~0_combout ),
	.cout());
defparam \E_cmp_result~0 .lut_mask = 16'h6996;
defparam \E_cmp_result~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_invert_arith_src_msb~0 (
	.dataa(\Equal0~8_combout ),
	.datab(\Equal62~0_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~0_combout ),
	.cout());
defparam \E_invert_arith_src_msb~0 .lut_mask = 16'hEFFE;
defparam \E_invert_arith_src_msb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_invert_arith_src_msb~1 (
	.dataa(\R_valid~q ),
	.datab(\E_invert_arith_src_msb~0_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_alu_subtract~8_combout ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~1_combout ),
	.cout());
defparam \E_invert_arith_src_msb~1 .lut_mask = 16'hEFFF;
defparam \E_invert_arith_src_msb~1 .sum_lutc_input = "datac";

dffeas E_invert_arith_src_msb(
	.clk(wire_pll7_clk_0),
	.d(\E_invert_arith_src_msb~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_invert_arith_src_msb~q ),
	.prn(vcc));
defparam E_invert_arith_src_msb.is_wysiwyg = "true";
defparam E_invert_arith_src_msb.power_up = "low";

cycloneive_lcell_comb \Add1~83 (
	.dataa(\E_alu_sub~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add1~83_combout ),
	.cout());
defparam \Add1~83 .lut_mask = 16'h9696;
defparam \Add1~83 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_arith_src1[31] (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(\E_src1[31]~q ),
	.cin(gnd),
	.combout(\E_arith_src1[31]~combout ),
	.cout());
defparam \E_arith_src1[31] .lut_mask = 16'h0FF0;
defparam \E_arith_src1[31] .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~84 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[30]~q ),
	.cin(gnd),
	.combout(\Add1~84_combout ),
	.cout());
defparam \Add1~84 .lut_mask = 16'h0FF0;
defparam \Add1~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[29]~q ),
	.cin(gnd),
	.combout(\Add1~85_combout ),
	.cout());
defparam \Add1~85 .lut_mask = 16'h0FF0;
defparam \Add1~85 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~86 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[28]~q ),
	.cin(gnd),
	.combout(\Add1~86_combout ),
	.cout());
defparam \Add1~86 .lut_mask = 16'h0FF0;
defparam \Add1~86 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~87 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[27]~q ),
	.cin(gnd),
	.combout(\Add1~87_combout ),
	.cout());
defparam \Add1~87 .lut_mask = 16'h0FF0;
defparam \Add1~87 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~98 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~97 ),
	.combout(\Add1~98_combout ),
	.cout());
defparam \Add1~98 .lut_mask = 16'h5A5A;
defparam \Add1~98 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_cmp_result~1 (
	.dataa(\E_cmp_result~0_combout ),
	.datab(\R_compare_op[1]~q ),
	.datac(\Add1~98_combout ),
	.datad(\R_compare_op[0]~q ),
	.cin(gnd),
	.combout(\E_cmp_result~1_combout ),
	.cout());
defparam \E_cmp_result~1 .lut_mask = 16'hEBBE;
defparam \E_cmp_result~1 .sum_lutc_input = "datac";

dffeas W_cmp_result(
	.clk(wire_pll7_clk_0),
	.d(\E_cmp_result~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_cmp_result~q ),
	.prn(vcc));
defparam W_cmp_result.is_wysiwyg = "true";
defparam W_cmp_result.power_up = "low";

cycloneive_lcell_comb \F_pc_sel_nxt~0 (
	.dataa(\R_ctrl_uncond_cti_non_br~q ),
	.datab(\R_ctrl_br_uncond~q ),
	.datac(\W_cmp_result~q ),
	.datad(\R_ctrl_br~q ),
	.cin(gnd),
	.combout(\F_pc_sel_nxt~0_combout ),
	.cout());
defparam \F_pc_sel_nxt~0 .lut_mask = 16'hFFFE;
defparam \F_pc_sel_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[24]~0 (
	.dataa(\R_ctrl_break~q ),
	.datab(\F_pc_plus_one[24]~48_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[24]~0_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[24]~0 .lut_mask = 16'hEFFF;
defparam \F_pc_no_crst_nxt[24]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[24]~1 (
	.dataa(\F_pc_no_crst_nxt[24]~0_combout ),
	.datab(\Add1~81_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[24]~1_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[24]~1 .lut_mask = 16'hFF7F;
defparam \F_pc_no_crst_nxt[24]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[23]~2 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\F_pc_plus_one[23]~46_combout ),
	.datac(\R_ctrl_break~q ),
	.datad(\F_pc_sel_nxt~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[23]~2_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[23]~2 .lut_mask = 16'hEFFF;
defparam \F_pc_no_crst_nxt[23]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[23]~3 (
	.dataa(\F_pc_no_crst_nxt[23]~2_combout ),
	.datab(\Add1~79_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[23]~3_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[23]~3 .lut_mask = 16'hFEFF;
defparam \F_pc_no_crst_nxt[23]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[22]~4 (
	.dataa(\Add1~77_combout ),
	.datab(\F_pc_plus_one[22]~44_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[22]~4_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[22]~4 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[22]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[21]~5 (
	.dataa(\Add1~75_combout ),
	.datab(\F_pc_plus_one[21]~42_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[21]~5_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[21]~5 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[21]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[20]~6 (
	.dataa(\Add1~73_combout ),
	.datab(\F_pc_plus_one[20]~40_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[20]~6_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[20]~6 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[20]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[19]~7 (
	.dataa(\Add1~71_combout ),
	.datab(\F_pc_plus_one[19]~38_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[19]~7_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[19]~7 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[19]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[18]~8 (
	.dataa(\Add1~69_combout ),
	.datab(\F_pc_plus_one[18]~36_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[18]~8_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[18]~8 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[18]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[17]~9 (
	.dataa(\Add1~67_combout ),
	.datab(\F_pc_plus_one[17]~34_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[17]~9_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[17]~9 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[17]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[16]~10 (
	.dataa(\Add1~65_combout ),
	.datab(\F_pc_plus_one[16]~32_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[16]~10_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[16]~10 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[16]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[15]~11 (
	.dataa(\Add1~63_combout ),
	.datab(\F_pc_plus_one[15]~30_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[15]~11_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[15]~11 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[15]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[14]~12 (
	.dataa(\Add1~61_combout ),
	.datab(\F_pc_plus_one[14]~28_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[14]~12_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[14]~12 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[14]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[13]~13 (
	.dataa(\Add1~59_combout ),
	.datab(\F_pc_plus_one[13]~26_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[13]~13_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[13]~13 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[13]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[12]~14 (
	.dataa(\Add1~57_combout ),
	.datab(\F_pc_plus_one[12]~24_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[12]~14_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[12]~14 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[12]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[11]~15 (
	.dataa(\Add1~55_combout ),
	.datab(\F_pc_plus_one[11]~22_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[11]~15_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[11]~15 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[11]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[10]~16 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(\F_pc_sel_nxt.10~0_combout ),
	.datac(\F_pc_plus_one[10]~20_combout ),
	.datad(\Add1~53_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[10]~16_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[10]~16 .lut_mask = 16'hFFF6;
defparam \F_pc_no_crst_nxt[10]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[10]~17 (
	.dataa(\R_ctrl_break~q ),
	.datab(\R_ctrl_exception~q ),
	.datac(\F_pc_no_crst_nxt[10]~16_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[10]~17_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[10]~17 .lut_mask = 16'hDFDF;
defparam \F_pc_no_crst_nxt[10]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[8]~18 (
	.dataa(\Add1~49_combout ),
	.datab(\F_pc_plus_one[8]~16_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[8]~18_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[8]~18 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[8]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[9]~19 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(\F_pc_sel_nxt.10~0_combout ),
	.datac(\F_pc_plus_one[9]~18_combout ),
	.datad(\Add1~51_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[9]~19_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[9]~19 .lut_mask = 16'hFFF6;
defparam \F_pc_no_crst_nxt[9]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[9]~20 (
	.dataa(\R_ctrl_break~q ),
	.datab(\R_ctrl_exception~q ),
	.datac(\F_pc_no_crst_nxt[9]~19_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[9]~20_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[9]~20 .lut_mask = 16'hFBFB;
defparam \F_pc_no_crst_nxt[9]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[0]~21 (
	.dataa(\Add1~13_combout ),
	.datab(\F_pc_plus_one[0]~0_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[0]~21_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[0]~21 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[0]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[1]~22 (
	.dataa(\Add1~15_combout ),
	.datab(\F_pc_plus_one[1]~2_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[1]~22_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[1]~22 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[1]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[2]~23 (
	.dataa(\Add1~17_combout ),
	.datab(\F_pc_plus_one[2]~4_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[2]~23_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[2]~23 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[2]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[3]~24 (
	.dataa(\F_pc_sel_nxt.10~0_combout ),
	.datab(\Add1~19_combout ),
	.datac(\F_pc_plus_one[3]~6_combout ),
	.datad(\F_pc_sel_nxt~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[3]~24_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[3]~24 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[3]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[4]~25 (
	.dataa(\Add1~21_combout ),
	.datab(\F_pc_plus_one[4]~8_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[4]~25_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[4]~25 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[4]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[5]~26 (
	.dataa(\Add1~43_combout ),
	.datab(\F_pc_plus_one[5]~10_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[5]~26_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[5]~26 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[5]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[6]~27 (
	.dataa(\Add1~45_combout ),
	.datab(\F_pc_plus_one[6]~12_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[6]~27_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[6]~27 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[6]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[7]~28 (
	.dataa(\Add1~47_combout ),
	.datab(\F_pc_plus_one[7]~14_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[7]~28_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[7]~28 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[7]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[10]~0 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[10]~0_combout ),
	.cout());
defparam \E_st_data[10]~0 .lut_mask = 16'hEFFE;
defparam \E_st_data[10]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[2]~2 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~11_combout ),
	.datac(\D_ctrl_mem8~1_combout ),
	.datad(\Add1~9_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[2]~2_combout ),
	.cout());
defparam \E_mem_byte_en[2]~2 .lut_mask = 16'hDEFF;
defparam \E_mem_byte_en[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[3]~3 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~11_combout ),
	.datac(\Add1~9_combout ),
	.datad(\D_ctrl_mem8~1_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[3]~3_combout ),
	.cout());
defparam \E_mem_byte_en[3]~3 .lut_mask = 16'hFDFE;
defparam \E_mem_byte_en[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \hbreak_enabled~0 (
	.dataa(\D_op_cmpge~0_combout ),
	.datab(\Equal62~9_combout ),
	.datac(hbreak_enabled1),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.cout());
defparam \hbreak_enabled~0 .lut_mask = 16'hFFF7;
defparam \hbreak_enabled~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[8]~1 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[8]~1_combout ),
	.cout());
defparam \E_st_data[8]~1 .lut_mask = 16'hEFFE;
defparam \E_st_data[8]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[9]~2 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[9]~2_combout ),
	.cout());
defparam \E_st_data[9]~2 .lut_mask = 16'hEFFE;
defparam \E_st_data[9]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[11]~3 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[11]~3_combout ),
	.cout());
defparam \E_st_data[11]~3 .lut_mask = 16'hEFFE;
defparam \E_st_data[11]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[12]~4 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[12]~4_combout ),
	.cout());
defparam \E_st_data[12]~4 .lut_mask = 16'hEFFE;
defparam \E_st_data[12]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[13]~5 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[13]~5_combout ),
	.cout());
defparam \E_st_data[13]~5 .lut_mask = 16'hEFFE;
defparam \E_st_data[13]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[14]~6 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[14]~6_combout ),
	.cout());
defparam \E_st_data[14]~6 .lut_mask = 16'hEFFE;
defparam \E_st_data[14]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[15]~7 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[15]~7_combout ),
	.cout());
defparam \E_st_data[15]~7 .lut_mask = 16'hEFFE;
defparam \E_st_data[15]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_byteenable[3]~0 (
	.dataa(\D_ctrl_mem8~0_combout ),
	.datab(\D_ctrl_mem16~0_combout ),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\d_byteenable[3]~0_combout ),
	.cout());
defparam \d_byteenable[3]~0 .lut_mask = 16'hEEFF;
defparam \d_byteenable[3]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[16]~8 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[16]~8_combout ),
	.cout());
defparam \E_st_data[16]~8 .lut_mask = 16'hAACC;
defparam \E_st_data[16]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[17]~9 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[17]~9_combout ),
	.cout());
defparam \E_st_data[17]~9 .lut_mask = 16'hAACC;
defparam \E_st_data[17]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[18]~10 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[18]~10_combout ),
	.cout());
defparam \E_st_data[18]~10 .lut_mask = 16'hAACC;
defparam \E_st_data[18]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[19]~11 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[19]~11_combout ),
	.cout());
defparam \E_st_data[19]~11 .lut_mask = 16'hAACC;
defparam \E_st_data[19]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[20]~12 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[20]~12_combout ),
	.cout());
defparam \E_st_data[20]~12 .lut_mask = 16'hAACC;
defparam \E_st_data[20]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[21]~13 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[21]~13_combout ),
	.cout());
defparam \E_st_data[21]~13 .lut_mask = 16'hAACC;
defparam \E_st_data[21]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[22]~14 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[22]~14_combout ),
	.cout());
defparam \E_st_data[22]~14 .lut_mask = 16'hAACC;
defparam \E_st_data[22]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[23]~15 (
	.dataa(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datab(\niosII_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[23]~15_combout ),
	.cout());
defparam \E_st_data[23]~15 .lut_mask = 16'hAACC;
defparam \E_st_data[23]~15 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_cpu_cpu_nios2_oci (
	wire_pll7_clk_0,
	sr_0,
	jtag_break,
	readdata_4,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	hbreak_enabled,
	WideOr1,
	rf_source_valid,
	uav_write,
	r_early_rst,
	address_nxt,
	oci_ienable_4,
	oci_ienable_3,
	oci_ienable_2,
	oci_ienable_1,
	oci_ienable_0,
	oci_single_step_mode,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	debugaccess_nxt,
	writedata_nxt,
	byteenable_nxt,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_14,
	readdata_15,
	readdata_10,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_6,
	readdata_21,
	readdata_30,
	readdata_29,
	readdata_28,
	readdata_27,
	readdata_26,
	readdata_25,
	readdata_24,
	readdata_23,
	readdata_22,
	readdata_20,
	readdata_19,
	readdata_18,
	readdata_17,
	readdata_31,
	resetrequest,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	sr_0;
output 	jtag_break;
output 	readdata_4;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
input 	saved_grant_0;
output 	waitrequest;
input 	mem_used_1;
input 	hbreak_enabled;
input 	WideOr1;
input 	rf_source_valid;
input 	uav_write;
input 	r_early_rst;
input 	[8:0] address_nxt;
output 	oci_ienable_4;
output 	oci_ienable_3;
output 	oci_ienable_2;
output 	oci_ienable_1;
output 	oci_ienable_0;
output 	oci_single_step_mode;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
input 	debugaccess_nxt;
input 	[31:0] writedata_nxt;
input 	[3:0] byteenable_nxt;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_5;
output 	readdata_14;
output 	readdata_15;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_6;
output 	readdata_21;
output 	readdata_30;
output 	readdata_29;
output 	readdata_28;
output 	readdata_27;
output 	readdata_26;
output 	readdata_25;
output 	readdata_24;
output 	readdata_23;
output 	readdata_22;
output 	readdata_20;
output 	readdata_19;
output 	readdata_18;
output 	readdata_17;
output 	readdata_31;
output 	resetrequest;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[0]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[1]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[3]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[4]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[25]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[26]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[5]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[29]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[11]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[12]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[9]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[8]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[18]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[0]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[1]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[0]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[36]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[37]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|ir[0]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|ir[1]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|enable_action_strobe~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[3]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ;
wire \the_niosII_cpu_cpu_nios2_oci_debug|monitor_ready~q ;
wire \write~q ;
wire \read~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[2]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[2]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[1]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[4]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[26]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[34]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[28]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[27]~q ;
wire \debugaccess~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|ociram_wr_en~0_combout ;
wire \writedata[0]~q ;
wire \address[1]~q ;
wire \address[2]~q ;
wire \address[3]~q ;
wire \address[4]~q ;
wire \address[5]~q ;
wire \address[6]~q ;
wire \address[7]~q ;
wire \byteenable[0]~q ;
wire \the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~0_combout ;
wire \the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ;
wire \the_niosII_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[25]~q ;
wire \write~0_combout ;
wire \write~1_combout ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[17]~q ;
wire \read~0_combout ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[21]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[20]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[3]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[2]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[5]~q ;
wire \writedata[1]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[29]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[30]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[31]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[32]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[33]~q ;
wire \writedata[4]~q ;
wire \writedata[3]~q ;
wire \writedata[2]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[19]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[18]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_debug|monitor_error~q ;
wire \the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ;
wire \the_niosII_cpu_cpu_nios2_oci_debug|monitor_go~q ;
wire \the_niosII_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[4]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[6]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[25]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[27]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[27]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[26]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[24]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[24]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[16]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[16]~q ;
wire \the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[23]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[20]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[20]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[19]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[19]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[23]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[5]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[7]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[28]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[28]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[29]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[30]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[30]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[31]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[31]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_debug|resetlatch~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[24]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[17]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[17]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[16]~q ;
wire \writedata[11]~q ;
wire \byteenable[1]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[13]~q ;
wire \writedata[13]~q ;
wire \writedata[16]~q ;
wire \byteenable[2]~q ;
wire \writedata[12]~q ;
wire \writedata[5]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[14]~q ;
wire \writedata[14]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[15]~q ;
wire \writedata[15]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[10]~q ;
wire \writedata[10]~q ;
wire \writedata[9]~q ;
wire \writedata[8]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[7]~q ;
wire \writedata[7]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[6]~q ;
wire \writedata[6]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[21]~q ;
wire \writedata[21]~q ;
wire \writedata[30]~q ;
wire \byteenable[3]~q ;
wire \writedata[29]~q ;
wire \writedata[28]~q ;
wire \writedata[27]~q ;
wire \writedata[26]~q ;
wire \writedata[25]~q ;
wire \writedata[24]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[23]~q ;
wire \writedata[23]~q ;
wire \the_niosII_cpu_cpu_nios2_ocimem|MonDReg[22]~q ;
wire \writedata[22]~q ;
wire \writedata[20]~q ;
wire \writedata[19]~q ;
wire \writedata[18]~q ;
wire \writedata[17]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[22]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[18]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[21]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[6]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[8]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[14]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[15]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[13]~q ;
wire \writedata[31]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[12]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[11]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[10]~q ;
wire \the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[9]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[22]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[7]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[23]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[15]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[8]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[13]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[14]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[12]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[11]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[10]~q ;
wire \the_niosII_cpu_cpu_nios2_oci_break|break_readreg[9]~q ;
wire \address[8]~q ;
wire \readdata~0_combout ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;
wire \readdata~3_combout ;
wire \readdata~4_combout ;
wire \readdata~5_combout ;
wire \readdata~6_combout ;
wire \readdata~7_combout ;
wire \readdata~8_combout ;
wire \address[0]~q ;
wire \readdata~9_combout ;
wire \readdata~10_combout ;
wire \readdata~11_combout ;
wire \readdata~12_combout ;
wire \readdata~13_combout ;
wire \readdata~14_combout ;
wire \readdata~15_combout ;
wire \readdata~16_combout ;
wire \readdata~17_combout ;
wire \readdata~18_combout ;
wire \readdata~19_combout ;
wire \readdata~20_combout ;
wire \readdata~21_combout ;
wire \readdata~22_combout ;
wire \readdata~23_combout ;
wire \readdata~24_combout ;
wire \readdata~25_combout ;
wire \readdata~26_combout ;
wire \readdata~27_combout ;
wire \readdata~28_combout ;
wire \readdata~29_combout ;
wire \readdata~30_combout ;
wire \readdata~31_combout ;
wire \readdata~32_combout ;
wire \readdata~33_combout ;
wire \readdata~34_combout ;
wire \readdata~35_combout ;
wire \readdata~36_combout ;
wire \readdata~37_combout ;


niosII_niosII_cpu_cpu_nios2_oci_break the_niosII_cpu_cpu_nios2_oci_break(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.break_readreg_0(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[1]~q ),
	.jdo_0(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_0(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|ir[0]~q ),
	.ir_1(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|ir[1]~q ),
	.enable_action_strobe(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.break_readreg_2(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[2]~q ),
	.jdo_1(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_25(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_17(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_21(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.break_readreg_3(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[3]~q ),
	.jdo_2(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_29(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_19(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.break_readreg_4(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_25(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_27(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_26(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_24(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_16(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_20(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[19]~q ),
	.jdo_23(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.break_readreg_5(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_7(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.break_readreg_28(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_29(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[31]~q ),
	.jdo_24(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.break_readreg_17(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[17]~q ),
	.jdo_16(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.jdo_22(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.break_readreg_18(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_21(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_6(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[6]~q ),
	.jdo_8(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_14(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_13(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_22(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_7(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_23(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_15(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_8(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_13(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[9]~q ));

niosII_niosII_cpu_cpu_nios2_oci_debug the_niosII_cpu_cpu_nios2_oci_debug(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.jtag_break1(jtag_break),
	.r_sync_rst(r_sync_rst),
	.take_action_ocimem_a(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.monitor_ready1(\the_niosII_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.jdo_34(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.writedata_0(\writedata[0]~q ),
	.take_action_ocireg(\the_niosII_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_25(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_21(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.take_action_ocimem_a1(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.writedata_1(\writedata[1]~q ),
	.jdo_19(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.monitor_error1(\the_niosII_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.monitor_go1(\the_niosII_cpu_cpu_nios2_oci_debug|monitor_go~q ),
	.resetrequest1(resetrequest),
	.jdo_23(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.resetlatch1(\the_niosII_cpu_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_24(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_22(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.state_1(state_1));

niosII_niosII_cpu_cpu_nios2_ocimem the_niosII_cpu_cpu_nios2_ocimem(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.MonDReg_0(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[0]~q ),
	.MonDReg_1(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[1]~q ),
	.q_a_0(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.MonDReg_3(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[3]~q ),
	.q_a_2(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.MonDReg_4(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_25(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_26(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[26]~q ),
	.q_a_11(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_12(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_5(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_14(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_10(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_8(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_7(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_21(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_30(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_29(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_28(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_27(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_26(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_25(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_24(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_23(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_22(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_20(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_18(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.MonDReg_5(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_29(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[29]~q ),
	.MonDReg_11(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_12(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[12]~q ),
	.q_a_31(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.MonDReg_9(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_8(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_18(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[18]~q ),
	.waitrequest1(waitrequest),
	.jdo_3(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.take_action_ocimem_b(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.take_no_action_ocimem_a(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.MonDReg_2(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[2]~q ),
	.jdo_4(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_34(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.take_action_ocimem_a(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_28(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.debugaccess(\debugaccess~q ),
	.ociram_wr_en(\the_niosII_cpu_cpu_nios2_ocimem|ociram_wr_en~0_combout ),
	.r_early_rst(r_early_rst),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.byteenable_0(\byteenable[0]~q ),
	.jdo_25(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_17(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_21(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_5(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_29(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_32(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_33(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[33]~q ),
	.writedata_4(\writedata[4]~q ),
	.writedata_3(\writedata[3]~q ),
	.writedata_2(\writedata[2]~q ),
	.jdo_19(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.jdo_6(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.MonDReg_27(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[27]~q ),
	.MonDReg_24(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[24]~q ),
	.MonDReg_16(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[16]~q ),
	.MonDReg_20(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[19]~q ),
	.jdo_23(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_7(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.MonDReg_28(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_30(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_31(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[31]~q ),
	.jdo_24(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.MonDReg_17(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[17]~q ),
	.jdo_16(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.writedata_11(\writedata[11]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.MonDReg_13(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[13]~q ),
	.writedata_13(\writedata[13]~q ),
	.writedata_16(\writedata[16]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.writedata_12(\writedata[12]~q ),
	.writedata_5(\writedata[5]~q ),
	.MonDReg_14(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[14]~q ),
	.writedata_14(\writedata[14]~q ),
	.MonDReg_15(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[15]~q ),
	.writedata_15(\writedata[15]~q ),
	.MonDReg_10(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[10]~q ),
	.writedata_10(\writedata[10]~q ),
	.writedata_9(\writedata[9]~q ),
	.writedata_8(\writedata[8]~q ),
	.MonDReg_7(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[7]~q ),
	.writedata_7(\writedata[7]~q ),
	.MonDReg_6(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[6]~q ),
	.writedata_6(\writedata[6]~q ),
	.MonDReg_21(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[21]~q ),
	.writedata_21(\writedata[21]~q ),
	.writedata_30(\writedata[30]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.writedata_29(\writedata[29]~q ),
	.writedata_28(\writedata[28]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_25(\writedata[25]~q ),
	.writedata_24(\writedata[24]~q ),
	.MonDReg_23(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[23]~q ),
	.writedata_23(\writedata[23]~q ),
	.MonDReg_22(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[22]~q ),
	.writedata_22(\writedata[22]~q ),
	.writedata_20(\writedata[20]~q ),
	.writedata_19(\writedata[19]~q ),
	.writedata_18(\writedata[18]~q ),
	.writedata_17(\writedata[17]~q ),
	.jdo_22(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_8(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_14(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_13(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.writedata_31(\writedata[31]~q ),
	.jdo_12(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[9]~q ));

niosII_niosII_cpu_cpu_nios2_avalon_reg the_niosII_cpu_cpu_nios2_avalon_reg(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.address_8(\address[8]~q ),
	.ociram_wr_en(\the_niosII_cpu_cpu_nios2_ocimem|ociram_wr_en~0_combout ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.Equal0(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~0_combout ),
	.Equal01(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.take_action_ocireg(\the_niosII_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.oci_ienable_4(oci_ienable_4),
	.oci_ienable_3(oci_ienable_3),
	.oci_ienable_2(oci_ienable_2),
	.oci_ienable_1(oci_ienable_1),
	.oci_ienable_0(oci_ienable_0),
	.oci_single_step_mode1(oci_single_step_mode),
	.writedata_1(\writedata[1]~q ),
	.writedata_4(\writedata[4]~q ),
	.writedata_3(\writedata[3]~q ),
	.writedata_2(\writedata[2]~q ),
	.Equal02(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.oci_reg_readdata(\the_niosII_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.oci_ienable_23(\the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[23]~q ));

niosII_niosII_cpu_cpu_debug_slave_wrapper the_niosII_cpu_cpu_debug_slave_wrapper(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.sr_0(sr_0),
	.MonDReg_0(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[0]~q ),
	.MonDReg_1(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[1]~q ),
	.MonDReg_3(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[3]~q ),
	.MonDReg_4(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_25(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_26(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_5(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_29(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[29]~q ),
	.MonDReg_11(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_12(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_9(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_8(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_18(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[18]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.break_readreg_0(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[1]~q ),
	.jdo_0(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_0(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|ir[0]~q ),
	.ir_1(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|ir[1]~q ),
	.enable_action_strobe(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.take_action_ocimem_b(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.take_action_ocimem_a(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.monitor_ready(\the_niosII_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.hbreak_enabled(hbreak_enabled),
	.break_readreg_2(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[2]~q ),
	.MonDReg_2(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[2]~q ),
	.jdo_1(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_34(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.take_action_ocimem_a1(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_28(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_25(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_17(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_21(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.take_action_ocimem_a2(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.break_readreg_3(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[3]~q ),
	.jdo_2(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_29(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_32(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_33(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_19(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.monitor_error(\the_niosII_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.break_readreg_4(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_25(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_27(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[27]~q ),
	.MonDReg_27(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[27]~q ),
	.break_readreg_26(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_24(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_16(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_20(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[19]~q ),
	.jdo_23(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.break_readreg_5(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_7(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.break_readreg_28(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[28]~q ),
	.MonDReg_28(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[28]~q ),
	.break_readreg_29(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[30]~q ),
	.MonDReg_30(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[30]~q ),
	.break_readreg_31(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[31]~q ),
	.MonDReg_31(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[31]~q ),
	.resetlatch(\the_niosII_cpu_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_24(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.break_readreg_17(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[17]~q ),
	.MonDReg_17(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[17]~q ),
	.jdo_16(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.MonDReg_13(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_15(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_10(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_7(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_6(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_21(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[21]~q ),
	.MonDReg_23(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_22(\the_niosII_cpu_cpu_nios2_ocimem|MonDReg[22]~q ),
	.jdo_22(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.break_readreg_18(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_21(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_6(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[6]~q ),
	.jdo_8(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_14(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_13(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_niosII_cpu_cpu_debug_slave_wrapper|the_niosII_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_22(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_7(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_23(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_15(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_8(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_13(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_niosII_cpu_cpu_nios2_oci_break|break_readreg[9]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

dffeas write(
	.clk(wire_pll7_clk_0),
	.d(\write~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(wire_pll7_clk_0),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas debugaccess(
	.clk(wire_pll7_clk_0),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \writedata[0] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \address[1] (
	.clk(wire_pll7_clk_0),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[2] (
	.clk(wire_pll7_clk_0),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[3] (
	.clk(wire_pll7_clk_0),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[4] (
	.clk(wire_pll7_clk_0),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \address[5] (
	.clk(wire_pll7_clk_0),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[6] (
	.clk(wire_pll7_clk_0),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[7] (
	.clk(wire_pll7_clk_0),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \byteenable[0] (
	.clk(wire_pll7_clk_0),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(uav_write),
	.datab(saved_grant_0),
	.datac(mem_used_1),
	.datad(\write~q ),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hEFFF;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~1 (
	.dataa(waitrequest),
	.datab(WideOr1),
	.datac(\write~0_combout ),
	.datad(\write~q ),
	.cin(gnd),
	.combout(\write~1_combout ),
	.cout());
defparam \write~1 .lut_mask = 16'hFFFE;
defparam \write~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(waitrequest),
	.datab(\read~q ),
	.datac(rf_source_valid),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hB8FF;
defparam \read~0 .sum_lutc_input = "datac";

dffeas \writedata[1] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[4] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[3] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \writedata[2] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[11] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \byteenable[1] (
	.clk(wire_pll7_clk_0),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[13] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[16] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \byteenable[2] (
	.clk(wire_pll7_clk_0),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[12] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[5] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[14] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[15] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[10] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[9] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[8] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[7] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[6] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[21] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[30] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \byteenable[3] (
	.clk(wire_pll7_clk_0),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[29] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \writedata[28] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[27] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[26] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[25] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[24] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \writedata[23] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[22] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \writedata[20] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \writedata[19] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \writedata[18] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[17] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[31] (
	.clk(wire_pll7_clk_0),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \readdata[4] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_cpu_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[0] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[11] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[13] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[16] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[12] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[5] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[14] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[10] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[9] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[8] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[7] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[6] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[21] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[30] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[29] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[28] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[27] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[26] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[25] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[24] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[23] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[22] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[20] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[19] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[18] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[17] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[31] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \address[8] (
	.clk(wire_pll7_clk_0),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cycloneive_lcell_comb \readdata~0 (
	.dataa(\address[8]~q ),
	.datab(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~0_combout ),
	.datac(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hFEFE;
defparam \readdata~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~1 (
	.dataa(\readdata~0_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.datac(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datad(oci_ienable_0),
	.cin(gnd),
	.combout(\readdata~1_combout ),
	.cout());
defparam \readdata~1 .lut_mask = 16'hACFF;
defparam \readdata~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~2 (
	.dataa(\readdata~1_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hEEFF;
defparam \readdata~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~3 (
	.dataa(\readdata~0_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.datac(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datad(oci_ienable_1),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hACFF;
defparam \readdata~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~4 (
	.dataa(\readdata~3_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hEEFF;
defparam \readdata~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~5 (
	.dataa(\readdata~0_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_oci_debug|monitor_go~q ),
	.datac(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datad(oci_ienable_2),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hACFF;
defparam \readdata~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~6 (
	.dataa(\readdata~5_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hEEFF;
defparam \readdata~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~7 (
	.dataa(\readdata~0_combout ),
	.datab(oci_single_step_mode),
	.datac(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datad(oci_ienable_3),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hACFF;
defparam \readdata~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~8 (
	.dataa(\readdata~7_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hEEFF;
defparam \readdata~8 .sum_lutc_input = "datac";

dffeas \address[0] (
	.clk(wire_pll7_clk_0),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

cycloneive_lcell_comb \readdata~9 (
	.dataa(\address[8]~q ),
	.datab(\the_niosII_cpu_cpu_nios2_avalon_reg|oci_ienable[23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata~9_combout ),
	.cout());
defparam \readdata~9 .lut_mask = 16'hEEEE;
defparam \readdata~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~10 (
	.dataa(\address[0]~q ),
	.datab(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~0_combout ),
	.datac(\the_niosII_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datad(\readdata~9_combout ),
	.cin(gnd),
	.combout(\readdata~10_combout ),
	.cout());
defparam \readdata~10 .lut_mask = 16'hFFFE;
defparam \readdata~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~11 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~11_combout ),
	.cout());
defparam \readdata~11 .lut_mask = 16'hEEFF;
defparam \readdata~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~12 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~12_combout ),
	.cout());
defparam \readdata~12 .lut_mask = 16'hEEFF;
defparam \readdata~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~13 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~13_combout ),
	.cout());
defparam \readdata~13 .lut_mask = 16'hEEFF;
defparam \readdata~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~14 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~14_combout ),
	.cout());
defparam \readdata~14 .lut_mask = 16'hEEFF;
defparam \readdata~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~15 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~15_combout ),
	.cout());
defparam \readdata~15 .lut_mask = 16'hEEFF;
defparam \readdata~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~16 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~16_combout ),
	.cout());
defparam \readdata~16 .lut_mask = 16'hEEFF;
defparam \readdata~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~17 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~17_combout ),
	.cout());
defparam \readdata~17 .lut_mask = 16'hEEFF;
defparam \readdata~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~18 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~18_combout ),
	.cout());
defparam \readdata~18 .lut_mask = 16'hEEFF;
defparam \readdata~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~19 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~19_combout ),
	.cout());
defparam \readdata~19 .lut_mask = 16'hEEFF;
defparam \readdata~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~20 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~20_combout ),
	.cout());
defparam \readdata~20 .lut_mask = 16'hEEFF;
defparam \readdata~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~21 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~21_combout ),
	.cout());
defparam \readdata~21 .lut_mask = 16'hEEFF;
defparam \readdata~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~22 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~22_combout ),
	.cout());
defparam \readdata~22 .lut_mask = 16'hEEFF;
defparam \readdata~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~23 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~23_combout ),
	.cout());
defparam \readdata~23 .lut_mask = 16'hEEFF;
defparam \readdata~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~24 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~24_combout ),
	.cout());
defparam \readdata~24 .lut_mask = 16'hEEFF;
defparam \readdata~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~25 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~25_combout ),
	.cout());
defparam \readdata~25 .lut_mask = 16'hEEFF;
defparam \readdata~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~26 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~26_combout ),
	.cout());
defparam \readdata~26 .lut_mask = 16'hEEFF;
defparam \readdata~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~27 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~27_combout ),
	.cout());
defparam \readdata~27 .lut_mask = 16'hEEFF;
defparam \readdata~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~28 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~28_combout ),
	.cout());
defparam \readdata~28 .lut_mask = 16'hEEFF;
defparam \readdata~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~29 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~29_combout ),
	.cout());
defparam \readdata~29 .lut_mask = 16'hEEFF;
defparam \readdata~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~30 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~30_combout ),
	.cout());
defparam \readdata~30 .lut_mask = 16'hEEFF;
defparam \readdata~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~31 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~31_combout ),
	.cout());
defparam \readdata~31 .lut_mask = 16'hEEFF;
defparam \readdata~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~32 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~32_combout ),
	.cout());
defparam \readdata~32 .lut_mask = 16'hEEFF;
defparam \readdata~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~33 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~33_combout ),
	.cout());
defparam \readdata~33 .lut_mask = 16'hEEFF;
defparam \readdata~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~34 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~34_combout ),
	.cout());
defparam \readdata~34 .lut_mask = 16'hEEFF;
defparam \readdata~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~35 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~35_combout ),
	.cout());
defparam \readdata~35 .lut_mask = 16'hEEFF;
defparam \readdata~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~36 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~36_combout ),
	.cout());
defparam \readdata~36 .lut_mask = 16'hEEFF;
defparam \readdata~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~37 (
	.dataa(\readdata~10_combout ),
	.datab(\the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~37_combout ),
	.cout());
defparam \readdata~37 .lut_mask = 16'hEEFF;
defparam \readdata~37 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_cpu_cpu_debug_slave_wrapper (
	wire_pll7_clk_0,
	sr_0,
	MonDReg_0,
	MonDReg_1,
	MonDReg_3,
	MonDReg_4,
	MonDReg_25,
	MonDReg_26,
	MonDReg_5,
	MonDReg_29,
	MonDReg_11,
	MonDReg_12,
	MonDReg_9,
	MonDReg_8,
	MonDReg_18,
	ir_out_0,
	ir_out_1,
	break_readreg_0,
	break_readreg_1,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_0,
	ir_1,
	enable_action_strobe,
	jdo_3,
	take_action_ocimem_b,
	take_action_ocimem_a,
	monitor_ready,
	hbreak_enabled,
	break_readreg_2,
	MonDReg_2,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_34,
	take_action_ocimem_a1,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_17,
	jdo_21,
	jdo_20,
	take_action_ocimem_a2,
	break_readreg_3,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_19,
	jdo_18,
	monitor_error,
	break_readreg_4,
	jdo_6,
	break_readreg_25,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	break_readreg_24,
	MonDReg_24,
	break_readreg_16,
	MonDReg_16,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	jdo_23,
	break_readreg_5,
	jdo_7,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	break_readreg_30,
	MonDReg_30,
	break_readreg_31,
	MonDReg_31,
	resetlatch,
	jdo_24,
	break_readreg_17,
	MonDReg_17,
	jdo_16,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_10,
	MonDReg_7,
	MonDReg_6,
	MonDReg_21,
	MonDReg_23,
	MonDReg_22,
	jdo_22,
	break_readreg_18,
	break_readreg_21,
	break_readreg_6,
	jdo_8,
	jdo_14,
	jdo_15,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_22,
	break_readreg_7,
	break_readreg_23,
	break_readreg_15,
	break_readreg_8,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	sr_0;
input 	MonDReg_0;
input 	MonDReg_1;
input 	MonDReg_3;
input 	MonDReg_4;
input 	MonDReg_25;
input 	MonDReg_26;
input 	MonDReg_5;
input 	MonDReg_29;
input 	MonDReg_11;
input 	MonDReg_12;
input 	MonDReg_9;
input 	MonDReg_8;
input 	MonDReg_18;
output 	ir_out_0;
output 	ir_out_1;
input 	break_readreg_0;
input 	break_readreg_1;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_0;
output 	ir_1;
output 	enable_action_strobe;
output 	jdo_3;
output 	take_action_ocimem_b;
output 	take_action_ocimem_a;
input 	monitor_ready;
input 	hbreak_enabled;
input 	break_readreg_2;
input 	MonDReg_2;
output 	jdo_1;
output 	jdo_4;
output 	jdo_26;
output 	jdo_34;
output 	take_action_ocimem_a1;
output 	jdo_28;
output 	jdo_27;
output 	jdo_25;
output 	jdo_17;
output 	jdo_21;
output 	jdo_20;
output 	take_action_ocimem_a2;
input 	break_readreg_3;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_19;
output 	jdo_18;
input 	monitor_error;
input 	break_readreg_4;
output 	jdo_6;
input 	break_readreg_25;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	jdo_23;
input 	break_readreg_5;
output 	jdo_7;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	break_readreg_30;
input 	MonDReg_30;
input 	break_readreg_31;
input 	MonDReg_31;
input 	resetlatch;
output 	jdo_24;
input 	break_readreg_17;
input 	MonDReg_17;
output 	jdo_16;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_10;
input 	MonDReg_7;
input 	MonDReg_6;
input 	MonDReg_21;
input 	MonDReg_23;
input 	MonDReg_22;
output 	jdo_22;
input 	break_readreg_18;
input 	break_readreg_21;
input 	break_readreg_6;
output 	jdo_8;
output 	jdo_14;
output 	jdo_15;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	break_readreg_22;
input 	break_readreg_7;
input 	break_readreg_23;
input 	break_readreg_15;
input 	break_readreg_8;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_niosII_cpu_cpu_debug_slave_tck|sr[35]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[31]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[7]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[15]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[1]~q ;
wire \niosII_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ;
wire \niosII_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[2]~q ;
wire \niosII_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[3]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[4]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[36]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[37]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[5]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[26]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[34]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[28]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[27]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[25]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[17]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[21]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[20]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[6]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[29]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[30]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[32]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[33]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[18]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[19]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[22]~q ;
wire \niosII_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[23]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[8]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[24]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[16]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[9]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[14]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[13]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[12]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[11]~q ;
wire \the_niosII_cpu_cpu_debug_slave_tck|sr[10]~q ;


niosII_niosII_cpu_cpu_debug_slave_sysclk the_niosII_cpu_cpu_debug_slave_sysclk(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.sr_0(sr_0),
	.sr_35(\the_niosII_cpu_cpu_debug_slave_tck|sr[35]~q ),
	.sr_31(\the_niosII_cpu_cpu_debug_slave_tck|sr[31]~q ),
	.sr_7(\the_niosII_cpu_cpu_debug_slave_tck|sr[7]~q ),
	.sr_15(\the_niosII_cpu_cpu_debug_slave_tck|sr[15]~q ),
	.sr_1(\the_niosII_cpu_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_niosII_cpu_cpu_debug_slave_tck|sr[2]~q ),
	.virtual_state_uir(\niosII_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.sr_3(\the_niosII_cpu_cpu_debug_slave_tck|sr[3]~q ),
	.jdo_0(jdo_0),
	.jdo_36(jdo_36),
	.jdo_37(jdo_37),
	.ir_0(ir_0),
	.ir_1(ir_1),
	.enable_action_strobe1(enable_action_strobe),
	.jdo_3(jdo_3),
	.take_action_ocimem_b1(take_action_ocimem_b),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.sr_4(\the_niosII_cpu_cpu_debug_slave_tck|sr[4]~q ),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_36(\the_niosII_cpu_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_niosII_cpu_cpu_debug_slave_tck|sr[37]~q ),
	.jdo_26(jdo_26),
	.jdo_34(jdo_34),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.jdo_28(jdo_28),
	.jdo_27(jdo_27),
	.jdo_25(jdo_25),
	.jdo_17(jdo_17),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.take_action_ocimem_a3(take_action_ocimem_a2),
	.sr_5(\the_niosII_cpu_cpu_debug_slave_tck|sr[5]~q ),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.sr_26(\the_niosII_cpu_cpu_debug_slave_tck|sr[26]~q ),
	.sr_34(\the_niosII_cpu_cpu_debug_slave_tck|sr[34]~q ),
	.sr_28(\the_niosII_cpu_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_niosII_cpu_cpu_debug_slave_tck|sr[27]~q ),
	.jdo_29(jdo_29),
	.jdo_30(jdo_30),
	.jdo_31(jdo_31),
	.jdo_32(jdo_32),
	.jdo_33(jdo_33),
	.sr_25(\the_niosII_cpu_cpu_debug_slave_tck|sr[25]~q ),
	.sr_17(\the_niosII_cpu_cpu_debug_slave_tck|sr[17]~q ),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.sr_21(\the_niosII_cpu_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_niosII_cpu_cpu_debug_slave_tck|sr[20]~q ),
	.sr_6(\the_niosII_cpu_cpu_debug_slave_tck|sr[6]~q ),
	.jdo_6(jdo_6),
	.sr_29(\the_niosII_cpu_cpu_debug_slave_tck|sr[29]~q ),
	.sr_30(\the_niosII_cpu_cpu_debug_slave_tck|sr[30]~q ),
	.sr_32(\the_niosII_cpu_cpu_debug_slave_tck|sr[32]~q ),
	.sr_33(\the_niosII_cpu_cpu_debug_slave_tck|sr[33]~q ),
	.sr_18(\the_niosII_cpu_cpu_debug_slave_tck|sr[18]~q ),
	.sr_19(\the_niosII_cpu_cpu_debug_slave_tck|sr[19]~q ),
	.sr_22(\the_niosII_cpu_cpu_debug_slave_tck|sr[22]~q ),
	.jdo_23(jdo_23),
	.jdo_7(jdo_7),
	.virtual_state_udr(\niosII_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.jdo_24(jdo_24),
	.jdo_16(jdo_16),
	.jdo_22(jdo_22),
	.sr_23(\the_niosII_cpu_cpu_debug_slave_tck|sr[23]~q ),
	.sr_8(\the_niosII_cpu_cpu_debug_slave_tck|sr[8]~q ),
	.jdo_8(jdo_8),
	.sr_24(\the_niosII_cpu_cpu_debug_slave_tck|sr[24]~q ),
	.sr_16(\the_niosII_cpu_cpu_debug_slave_tck|sr[16]~q ),
	.jdo_14(jdo_14),
	.jdo_15(jdo_15),
	.jdo_13(jdo_13),
	.jdo_12(jdo_12),
	.jdo_11(jdo_11),
	.jdo_10(jdo_10),
	.jdo_9(jdo_9),
	.sr_9(\the_niosII_cpu_cpu_debug_slave_tck|sr[9]~q ),
	.sr_14(\the_niosII_cpu_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_niosII_cpu_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_niosII_cpu_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_niosII_cpu_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_niosII_cpu_cpu_debug_slave_tck|sr[10]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}));

niosII_niosII_cpu_cpu_debug_slave_tck the_niosII_cpu_cpu_debug_slave_tck(
	.sr_0(sr_0),
	.MonDReg_0(MonDReg_0),
	.MonDReg_1(MonDReg_1),
	.sr_35(\the_niosII_cpu_cpu_debug_slave_tck|sr[35]~q ),
	.MonDReg_3(MonDReg_3),
	.MonDReg_4(MonDReg_4),
	.MonDReg_25(MonDReg_25),
	.MonDReg_26(MonDReg_26),
	.sr_31(\the_niosII_cpu_cpu_debug_slave_tck|sr[31]~q ),
	.sr_7(\the_niosII_cpu_cpu_debug_slave_tck|sr[7]~q ),
	.MonDReg_5(MonDReg_5),
	.MonDReg_29(MonDReg_29),
	.MonDReg_11(MonDReg_11),
	.MonDReg_12(MonDReg_12),
	.MonDReg_9(MonDReg_9),
	.MonDReg_8(MonDReg_8),
	.MonDReg_18(MonDReg_18),
	.sr_15(\the_niosII_cpu_cpu_debug_slave_tck|sr[15]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.sr_1(\the_niosII_cpu_cpu_debug_slave_tck|sr[1]~q ),
	.virtual_state_cdr(\niosII_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\niosII_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.sr_2(\the_niosII_cpu_cpu_debug_slave_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.virtual_state_uir(\niosII_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.sr_3(\the_niosII_cpu_cpu_debug_slave_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.monitor_ready(monitor_ready),
	.hbreak_enabled(hbreak_enabled),
	.sr_4(\the_niosII_cpu_cpu_debug_slave_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.MonDReg_2(MonDReg_2),
	.sr_36(\the_niosII_cpu_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_niosII_cpu_cpu_debug_slave_tck|sr[37]~q ),
	.sr_5(\the_niosII_cpu_cpu_debug_slave_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.sr_26(\the_niosII_cpu_cpu_debug_slave_tck|sr[26]~q ),
	.sr_34(\the_niosII_cpu_cpu_debug_slave_tck|sr[34]~q ),
	.sr_28(\the_niosII_cpu_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_niosII_cpu_cpu_debug_slave_tck|sr[27]~q ),
	.sr_25(\the_niosII_cpu_cpu_debug_slave_tck|sr[25]~q ),
	.sr_17(\the_niosII_cpu_cpu_debug_slave_tck|sr[17]~q ),
	.sr_21(\the_niosII_cpu_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_niosII_cpu_cpu_debug_slave_tck|sr[20]~q ),
	.monitor_error(monitor_error),
	.sr_6(\the_niosII_cpu_cpu_debug_slave_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.break_readreg_25(break_readreg_25),
	.sr_29(\the_niosII_cpu_cpu_debug_slave_tck|sr[29]~q ),
	.break_readreg_27(break_readreg_27),
	.MonDReg_27(MonDReg_27),
	.break_readreg_26(break_readreg_26),
	.sr_30(\the_niosII_cpu_cpu_debug_slave_tck|sr[30]~q ),
	.sr_32(\the_niosII_cpu_cpu_debug_slave_tck|sr[32]~q ),
	.sr_33(\the_niosII_cpu_cpu_debug_slave_tck|sr[33]~q ),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.sr_18(\the_niosII_cpu_cpu_debug_slave_tck|sr[18]~q ),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.sr_19(\the_niosII_cpu_cpu_debug_slave_tck|sr[19]~q ),
	.sr_22(\the_niosII_cpu_cpu_debug_slave_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.break_readreg_5(break_readreg_5),
	.break_readreg_28(break_readreg_28),
	.MonDReg_28(MonDReg_28),
	.break_readreg_29(break_readreg_29),
	.break_readreg_30(break_readreg_30),
	.MonDReg_30(MonDReg_30),
	.break_readreg_31(break_readreg_31),
	.MonDReg_31(MonDReg_31),
	.resetlatch(resetlatch),
	.break_readreg_17(break_readreg_17),
	.MonDReg_17(MonDReg_17),
	.MonDReg_13(MonDReg_13),
	.MonDReg_14(MonDReg_14),
	.MonDReg_15(MonDReg_15),
	.MonDReg_10(MonDReg_10),
	.MonDReg_7(MonDReg_7),
	.MonDReg_6(MonDReg_6),
	.MonDReg_21(MonDReg_21),
	.MonDReg_23(MonDReg_23),
	.MonDReg_22(MonDReg_22),
	.break_readreg_18(break_readreg_18),
	.sr_23(\the_niosII_cpu_cpu_debug_slave_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.break_readreg_6(break_readreg_6),
	.sr_8(\the_niosII_cpu_cpu_debug_slave_tck|sr[8]~q ),
	.sr_24(\the_niosII_cpu_cpu_debug_slave_tck|sr[24]~q ),
	.sr_16(\the_niosII_cpu_cpu_debug_slave_tck|sr[16]~q ),
	.break_readreg_22(break_readreg_22),
	.sr_9(\the_niosII_cpu_cpu_debug_slave_tck|sr[9]~q ),
	.break_readreg_7(break_readreg_7),
	.break_readreg_23(break_readreg_23),
	.break_readreg_15(break_readreg_15),
	.sr_14(\the_niosII_cpu_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_niosII_cpu_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_niosII_cpu_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_niosII_cpu_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_niosII_cpu_cpu_debug_slave_tck|sr[10]~q ),
	.break_readreg_8(break_readreg_8),
	.break_readreg_13(break_readreg_13),
	.break_readreg_14(break_readreg_14),
	.break_readreg_12(break_readreg_12),
	.break_readreg_11(break_readreg_11),
	.break_readreg_10(break_readreg_10),
	.break_readreg_9(break_readreg_9),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

niosII_sld_virtual_jtag_basic_1 niosII_cpu_cpu_debug_slave_phy(
	.virtual_state_cdr1(\niosII_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\niosII_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir(\niosII_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.virtual_state_udr(\niosII_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

endmodule

module niosII_niosII_cpu_cpu_debug_slave_sysclk (
	wire_pll7_clk_0,
	sr_0,
	sr_35,
	sr_31,
	sr_7,
	sr_15,
	sr_1,
	sr_2,
	virtual_state_uir,
	sr_3,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_0,
	ir_1,
	enable_action_strobe1,
	jdo_3,
	take_action_ocimem_b1,
	take_action_ocimem_a1,
	sr_4,
	jdo_1,
	jdo_4,
	sr_36,
	sr_37,
	jdo_26,
	jdo_34,
	take_action_ocimem_a2,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_17,
	jdo_21,
	jdo_20,
	take_action_ocimem_a3,
	sr_5,
	jdo_2,
	jdo_5,
	sr_26,
	sr_34,
	sr_28,
	sr_27,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	sr_25,
	sr_17,
	jdo_19,
	jdo_18,
	sr_21,
	sr_20,
	sr_6,
	jdo_6,
	sr_29,
	sr_30,
	sr_32,
	sr_33,
	sr_18,
	sr_19,
	sr_22,
	jdo_23,
	jdo_7,
	virtual_state_udr,
	jdo_24,
	jdo_16,
	jdo_22,
	sr_23,
	sr_8,
	jdo_8,
	sr_24,
	sr_16,
	jdo_14,
	jdo_15,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	sr_9,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	ir_in)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	sr_0;
input 	sr_35;
input 	sr_31;
input 	sr_7;
input 	sr_15;
input 	sr_1;
input 	sr_2;
input 	virtual_state_uir;
input 	sr_3;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_0;
output 	ir_1;
output 	enable_action_strobe1;
output 	jdo_3;
output 	take_action_ocimem_b1;
output 	take_action_ocimem_a1;
input 	sr_4;
output 	jdo_1;
output 	jdo_4;
input 	sr_36;
input 	sr_37;
output 	jdo_26;
output 	jdo_34;
output 	take_action_ocimem_a2;
output 	jdo_28;
output 	jdo_27;
output 	jdo_25;
output 	jdo_17;
output 	jdo_21;
output 	jdo_20;
output 	take_action_ocimem_a3;
input 	sr_5;
output 	jdo_2;
output 	jdo_5;
input 	sr_26;
input 	sr_34;
input 	sr_28;
input 	sr_27;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
input 	sr_25;
input 	sr_17;
output 	jdo_19;
output 	jdo_18;
input 	sr_21;
input 	sr_20;
input 	sr_6;
output 	jdo_6;
input 	sr_29;
input 	sr_30;
input 	sr_32;
input 	sr_33;
input 	sr_18;
input 	sr_19;
input 	sr_22;
output 	jdo_23;
output 	jdo_7;
input 	virtual_state_udr;
output 	jdo_24;
output 	jdo_16;
output 	jdo_22;
input 	sr_23;
input 	sr_8;
output 	jdo_8;
input 	sr_24;
input 	sr_16;
output 	jdo_14;
output 	jdo_15;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	sr_9;
input 	sr_14;
input 	sr_13;
input 	sr_12;
input 	sr_11;
input 	sr_10;
input 	[1:0] ir_in;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;
wire \jdo[35]~q ;


niosII_altera_std_synchronizer_2 the_altera_std_synchronizer3(
	.clk(wire_pll7_clk_0),
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr));

niosII_altera_std_synchronizer_3 the_altera_std_synchronizer4(
	.clk(wire_pll7_clk_0),
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ));

dffeas \jdo[0] (
	.clk(wire_pll7_clk_0),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[36] (
	.clk(wire_pll7_clk_0),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

dffeas \jdo[37] (
	.clk(wire_pll7_clk_0),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \ir[0] (
	.clk(wire_pll7_clk_0),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_0),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

dffeas \ir[1] (
	.clk(wire_pll7_clk_0),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_1),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas enable_action_strobe(
	.clk(wire_pll7_clk_0),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_action_strobe1),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

dffeas \jdo[3] (
	.clk(wire_pll7_clk_0),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

cycloneive_lcell_comb take_action_ocimem_b(
	.dataa(enable_action_strobe1),
	.datab(\jdo[35]~q ),
	.datac(ir_1),
	.datad(ir_0),
	.cin(gnd),
	.combout(take_action_ocimem_b1),
	.cout());
defparam take_action_ocimem_b.lut_mask = 16'hEFFF;
defparam take_action_ocimem_b.sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_ocimem_a~0 (
	.dataa(enable_action_strobe1),
	.datab(ir_1),
	.datac(ir_0),
	.datad(\jdo[35]~q ),
	.cin(gnd),
	.combout(take_action_ocimem_a1),
	.cout());
defparam \take_action_ocimem_a~0 .lut_mask = 16'hFFFD;
defparam \take_action_ocimem_a~0 .sum_lutc_input = "datac";

dffeas \jdo[1] (
	.clk(wire_pll7_clk_0),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(wire_pll7_clk_0),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[26] (
	.clk(wire_pll7_clk_0),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[34] (
	.clk(wire_pll7_clk_0),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

cycloneive_lcell_comb \take_action_ocimem_a~1 (
	.dataa(enable_action_strobe1),
	.datab(gnd),
	.datac(ir_1),
	.datad(ir_0),
	.cin(gnd),
	.combout(take_action_ocimem_a2),
	.cout());
defparam \take_action_ocimem_a~1 .lut_mask = 16'hAFFF;
defparam \take_action_ocimem_a~1 .sum_lutc_input = "datac";

dffeas \jdo[28] (
	.clk(wire_pll7_clk_0),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[27] (
	.clk(wire_pll7_clk_0),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[25] (
	.clk(wire_pll7_clk_0),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[17] (
	.clk(wire_pll7_clk_0),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

dffeas \jdo[21] (
	.clk(wire_pll7_clk_0),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(wire_pll7_clk_0),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

cycloneive_lcell_comb take_action_ocimem_a(
	.dataa(take_action_ocimem_a1),
	.datab(jdo_34),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(take_action_ocimem_a3),
	.cout());
defparam take_action_ocimem_a.lut_mask = 16'hDDDD;
defparam take_action_ocimem_a.sum_lutc_input = "datac";

dffeas \jdo[2] (
	.clk(wire_pll7_clk_0),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(wire_pll7_clk_0),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[29] (
	.clk(wire_pll7_clk_0),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[30] (
	.clk(wire_pll7_clk_0),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[31] (
	.clk(wire_pll7_clk_0),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[32] (
	.clk(wire_pll7_clk_0),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[33] (
	.clk(wire_pll7_clk_0),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[19] (
	.clk(wire_pll7_clk_0),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(wire_pll7_clk_0),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[6] (
	.clk(wire_pll7_clk_0),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[23] (
	.clk(wire_pll7_clk_0),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[7] (
	.clk(wire_pll7_clk_0),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[24] (
	.clk(wire_pll7_clk_0),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[16] (
	.clk(wire_pll7_clk_0),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[22] (
	.clk(wire_pll7_clk_0),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[8] (
	.clk(wire_pll7_clk_0),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[14] (
	.clk(wire_pll7_clk_0),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[15] (
	.clk(wire_pll7_clk_0),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[13] (
	.clk(wire_pll7_clk_0),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[12] (
	.clk(wire_pll7_clk_0),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas \jdo[11] (
	.clk(wire_pll7_clk_0),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[10] (
	.clk(wire_pll7_clk_0),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[9] (
	.clk(wire_pll7_clk_0),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas sync2_udr(
	.clk(wire_pll7_clk_0),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cycloneive_lcell_comb \update_jdo_strobe~0 (
	.dataa(\the_altera_std_synchronizer3|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_udr~q ),
	.cin(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.cout());
defparam \update_jdo_strobe~0 .lut_mask = 16'hAAFF;
defparam \update_jdo_strobe~0 .sum_lutc_input = "datac";

dffeas update_jdo_strobe(
	.clk(wire_pll7_clk_0),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(wire_pll7_clk_0),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cycloneive_lcell_comb \jxuir~0 (
	.dataa(\the_altera_std_synchronizer4|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_uir~q ),
	.cin(gnd),
	.combout(\jxuir~0_combout ),
	.cout());
defparam \jxuir~0 .lut_mask = 16'hAAFF;
defparam \jxuir~0 .sum_lutc_input = "datac";

dffeas jxuir(
	.clk(wire_pll7_clk_0),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

dffeas \jdo[35] (
	.clk(wire_pll7_clk_0),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(\jdo[35]~q ),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_2 (
	clk,
	dreg_0,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	dreg_0;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_3 (
	clk,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_niosII_cpu_cpu_debug_slave_tck (
	sr_0,
	MonDReg_0,
	MonDReg_1,
	sr_35,
	MonDReg_3,
	MonDReg_4,
	MonDReg_25,
	MonDReg_26,
	sr_31,
	sr_7,
	MonDReg_5,
	MonDReg_29,
	MonDReg_11,
	MonDReg_12,
	MonDReg_9,
	MonDReg_8,
	MonDReg_18,
	sr_15,
	ir_out_0,
	ir_out_1,
	sr_1,
	virtual_state_cdr,
	virtual_state_sdr,
	sr_2,
	break_readreg_0,
	virtual_state_uir,
	sr_3,
	break_readreg_1,
	monitor_ready,
	hbreak_enabled,
	sr_4,
	break_readreg_2,
	MonDReg_2,
	sr_36,
	sr_37,
	sr_5,
	break_readreg_3,
	sr_26,
	sr_34,
	sr_28,
	sr_27,
	sr_25,
	sr_17,
	sr_21,
	sr_20,
	monitor_error,
	sr_6,
	break_readreg_4,
	break_readreg_25,
	sr_29,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	sr_30,
	sr_32,
	sr_33,
	break_readreg_24,
	MonDReg_24,
	sr_18,
	break_readreg_16,
	MonDReg_16,
	sr_19,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	break_readreg_5,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	break_readreg_30,
	MonDReg_30,
	break_readreg_31,
	MonDReg_31,
	resetlatch,
	break_readreg_17,
	MonDReg_17,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_10,
	MonDReg_7,
	MonDReg_6,
	MonDReg_21,
	MonDReg_23,
	MonDReg_22,
	break_readreg_18,
	sr_23,
	break_readreg_21,
	break_readreg_6,
	sr_8,
	sr_24,
	sr_16,
	break_readreg_22,
	sr_9,
	break_readreg_7,
	break_readreg_23,
	break_readreg_15,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	break_readreg_8,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
input 	MonDReg_0;
input 	MonDReg_1;
output 	sr_35;
input 	MonDReg_3;
input 	MonDReg_4;
input 	MonDReg_25;
input 	MonDReg_26;
output 	sr_31;
output 	sr_7;
input 	MonDReg_5;
input 	MonDReg_29;
input 	MonDReg_11;
input 	MonDReg_12;
input 	MonDReg_9;
input 	MonDReg_8;
input 	MonDReg_18;
output 	sr_15;
output 	ir_out_0;
output 	ir_out_1;
output 	sr_1;
input 	virtual_state_cdr;
input 	virtual_state_sdr;
output 	sr_2;
input 	break_readreg_0;
input 	virtual_state_uir;
output 	sr_3;
input 	break_readreg_1;
input 	monitor_ready;
input 	hbreak_enabled;
output 	sr_4;
input 	break_readreg_2;
input 	MonDReg_2;
output 	sr_36;
output 	sr_37;
output 	sr_5;
input 	break_readreg_3;
output 	sr_26;
output 	sr_34;
output 	sr_28;
output 	sr_27;
output 	sr_25;
output 	sr_17;
output 	sr_21;
output 	sr_20;
input 	monitor_error;
output 	sr_6;
input 	break_readreg_4;
input 	break_readreg_25;
output 	sr_29;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
output 	sr_30;
output 	sr_32;
output 	sr_33;
input 	break_readreg_24;
input 	MonDReg_24;
output 	sr_18;
input 	break_readreg_16;
input 	MonDReg_16;
output 	sr_19;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	break_readreg_5;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	break_readreg_30;
input 	MonDReg_30;
input 	break_readreg_31;
input 	MonDReg_31;
input 	resetlatch;
input 	break_readreg_17;
input 	MonDReg_17;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_10;
input 	MonDReg_7;
input 	MonDReg_6;
input 	MonDReg_21;
input 	MonDReg_23;
input 	MonDReg_22;
input 	break_readreg_18;
output 	sr_23;
input 	break_readreg_21;
input 	break_readreg_6;
output 	sr_8;
output 	sr_24;
output 	sr_16;
input 	break_readreg_22;
output 	sr_9;
input 	break_readreg_7;
input 	break_readreg_23;
input 	break_readreg_15;
output 	sr_14;
output 	sr_13;
output 	sr_12;
output 	sr_11;
output 	sr_10;
input 	break_readreg_8;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \DRsize.000~q ;
wire \sr[0]~5_combout ;
wire \Mux37~0_combout ;
wire \sr~10_combout ;
wire \DRsize.100~q ;
wire \sr[35]~6_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr[31]~51_combout ;
wire \sr[31]~7_combout ;
wire \Mux30~0_combout ;
wire \sr[7]~8_combout ;
wire \sr[33]~83_combout ;
wire \DRsize.010~q ;
wire \sr[15]~9_combout ;
wire \sr~73_combout ;
wire \sr~74_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr[10]~13_combout ;
wire \sr~14_combout ;
wire \sr~15_combout ;
wire \sr~16_combout ;
wire \sr~17_combout ;
wire \sr~18_combout ;
wire \sr~19_combout ;
wire \sr~20_combout ;
wire \sr[37]~21_combout ;
wire \sr~22_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr~29_combout ;
wire \sr~30_combout ;
wire \sr[33]~31_combout ;
wire \sr~32_combout ;
wire \sr~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~36_combout ;
wire \sr~37_combout ;
wire \sr~38_combout ;
wire \sr~39_combout ;
wire \sr~40_combout ;
wire \sr~41_combout ;
wire \sr~42_combout ;
wire \sr~43_combout ;
wire \sr~44_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~48_combout ;
wire \sr~49_combout ;
wire \sr~50_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~55_combout ;
wire \sr~56_combout ;
wire \sr~57_combout ;
wire \sr~58_combout ;
wire \sr~59_combout ;
wire \sr~60_combout ;
wire \sr~61_combout ;
wire \sr~62_combout ;
wire \sr~63_combout ;
wire \sr~64_combout ;
wire \sr~65_combout ;
wire \sr~66_combout ;
wire \sr~67_combout ;
wire \sr~68_combout ;
wire \sr~69_combout ;
wire \sr~70_combout ;
wire \sr~71_combout ;
wire \sr~72_combout ;
wire \sr~75_combout ;
wire \sr~76_combout ;
wire \sr~77_combout ;
wire \sr~78_combout ;
wire \sr~79_combout ;
wire \sr~80_combout ;
wire \sr~81_combout ;
wire \sr~82_combout ;


niosII_altera_std_synchronizer_5 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

niosII_altera_std_synchronizer_4 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr[0]~5_combout ),
	.asdata(\sr~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr[35]~6_combout ),
	.asdata(\sr~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr[31]~7_combout ),
	.asdata(sr_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr[7]~8_combout ),
	.asdata(sr_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr[15]~9_combout ),
	.asdata(\sr~74_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~21_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~21_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~31_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[10]~13_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cycloneive_lcell_comb \sr[0]~5 (
	.dataa(altera_internal_jtag1),
	.datab(sr_1),
	.datac(gnd),
	.datad(\DRsize.000~q ),
	.cin(gnd),
	.combout(\sr[0]~5_combout ),
	.cout());
defparam \sr[0]~5 .lut_mask = 16'hAACC;
defparam \sr[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux37~0 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
defparam \Mux37~0 .lut_mask = 16'h7777;
defparam \Mux37~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~10 (
	.dataa(sr_0),
	.datab(virtual_state_cdr),
	.datac(\the_altera_std_synchronizer2|dreg[0]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~10_combout ),
	.cout());
defparam \sr~10 .lut_mask = 16'hFFB8;
defparam \sr~10 .sum_lutc_input = "datac";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cycloneive_lcell_comb \sr[35]~6 (
	.dataa(sr_36),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.100~q ),
	.cin(gnd),
	.combout(\sr[35]~6_combout ),
	.cout());
defparam \sr[35]~6 .lut_mask = 16'hAACC;
defparam \sr[35]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~23 (
	.dataa(irf_reg_1_2),
	.datab(state_3),
	.datac(splitter_nodes_receive_1_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~23_combout ),
	.cout());
defparam \sr~23 .lut_mask = 16'hFDFF;
defparam \sr~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~24 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(\the_altera_std_synchronizer1|dreg[0]~q ),
	.datad(\sr~23_combout ),
	.cin(gnd),
	.combout(\sr~24_combout ),
	.cout());
defparam \sr~24 .lut_mask = 16'hFFD8;
defparam \sr~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~25 (
	.dataa(sr_35),
	.datab(virtual_state_cdr),
	.datac(\sr~23_combout ),
	.datad(\sr~24_combout ),
	.cin(gnd),
	.combout(\sr~25_combout ),
	.cout());
defparam \sr~25 .lut_mask = 16'hFFFE;
defparam \sr~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[31]~51 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(break_readreg_30),
	.datad(MonDReg_30),
	.cin(gnd),
	.combout(\sr[31]~51_combout ),
	.cout());
defparam \sr[31]~51 .lut_mask = 16'hFFF6;
defparam \sr[31]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[31]~7 (
	.dataa(sr_31),
	.datab(virtual_state_cdr),
	.datac(irf_reg_0_2),
	.datad(\sr[31]~51_combout ),
	.cin(gnd),
	.combout(\sr[31]~7_combout ),
	.cout());
defparam \sr[31]~7 .lut_mask = 16'hBF8F;
defparam \sr[31]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux30~0 (
	.dataa(break_readreg_6),
	.datab(MonDReg_6),
	.datac(irf_reg_1_2),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
defparam \Mux30~0 .lut_mask = 16'hACFF;
defparam \Mux30~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[7]~8 (
	.dataa(\Mux30~0_combout ),
	.datab(sr_7),
	.datac(gnd),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\sr[7]~8_combout ),
	.cout());
defparam \sr[7]~8 .lut_mask = 16'hAACC;
defparam \sr[7]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[33]~83 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sr[33]~83_combout ),
	.cout());
defparam \sr[33]~83 .lut_mask = 16'hEEEE;
defparam \sr[33]~83 .sum_lutc_input = "datac";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[33]~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cycloneive_lcell_comb \sr[15]~9 (
	.dataa(sr_16),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.010~q ),
	.cin(gnd),
	.combout(\sr[15]~9_combout ),
	.cout());
defparam \sr[15]~9 .lut_mask = 16'hAACC;
defparam \sr[15]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~73 (
	.dataa(break_readreg_14),
	.datab(MonDReg_14),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~73_combout ),
	.cout());
defparam \sr~73 .lut_mask = 16'hAACC;
defparam \sr~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~74 (
	.dataa(sr_15),
	.datab(virtual_state_cdr),
	.datac(\sr~73_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~74_combout ),
	.cout());
defparam \sr~74 .lut_mask = 16'hB8FF;
defparam \sr~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~11 (
	.dataa(break_readreg_0),
	.datab(MonDReg_0),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~11_combout ),
	.cout());
defparam \sr~11 .lut_mask = 16'hAACC;
defparam \sr~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~12 (
	.dataa(sr_2),
	.datab(virtual_state_sdr),
	.datac(\sr~11_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~12_combout ),
	.cout());
defparam \sr~12 .lut_mask = 16'hB8FF;
defparam \sr~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[10]~13 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr[10]~13_combout ),
	.cout());
defparam \sr[10]~13 .lut_mask = 16'hFEFF;
defparam \sr[10]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~14 (
	.dataa(break_readreg_1),
	.datab(MonDReg_1),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~14_combout ),
	.cout());
defparam \sr~14 .lut_mask = 16'hAACC;
defparam \sr~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~15 (
	.dataa(sr_3),
	.datab(virtual_state_sdr),
	.datac(\sr~14_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~15_combout ),
	.cout());
defparam \sr~15 .lut_mask = 16'hB8FF;
defparam \sr~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~16 (
	.dataa(break_readreg_2),
	.datab(MonDReg_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~16_combout ),
	.cout());
defparam \sr~16 .lut_mask = 16'hAACC;
defparam \sr~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~17 (
	.dataa(sr_4),
	.datab(virtual_state_sdr),
	.datac(\sr~16_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~17_combout ),
	.cout());
defparam \sr~17 .lut_mask = 16'hB8FF;
defparam \sr~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~18 (
	.dataa(break_readreg_3),
	.datab(MonDReg_3),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~18_combout ),
	.cout());
defparam \sr~18 .lut_mask = 16'hAACC;
defparam \sr~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~19 (
	.dataa(sr_5),
	.datab(virtual_state_sdr),
	.datac(\sr~18_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~19_combout ),
	.cout());
defparam \sr~19 .lut_mask = 16'hB8FF;
defparam \sr~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~20 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(sr_37),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~20_combout ),
	.cout());
defparam \sr~20 .lut_mask = 16'hFEFF;
defparam \sr~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[37]~21 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[37]~21_combout ),
	.cout());
defparam \sr[37]~21 .lut_mask = 16'hFF7D;
defparam \sr[37]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~22 (
	.dataa(altera_internal_jtag1),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~22_combout ),
	.cout());
defparam \sr~22 .lut_mask = 16'hFEFF;
defparam \sr~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~26 (
	.dataa(break_readreg_4),
	.datab(MonDReg_4),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~26_combout ),
	.cout());
defparam \sr~26 .lut_mask = 16'hAACC;
defparam \sr~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~27 (
	.dataa(sr_6),
	.datab(virtual_state_sdr),
	.datac(\sr~26_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~27_combout ),
	.cout());
defparam \sr~27 .lut_mask = 16'hB8FF;
defparam \sr~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~28 (
	.dataa(break_readreg_25),
	.datab(MonDReg_25),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~28_combout ),
	.cout());
defparam \sr~28 .lut_mask = 16'hAACC;
defparam \sr~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~29 (
	.dataa(virtual_state_sdr),
	.datab(irf_reg_0_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~29_combout ),
	.cout());
defparam \sr~29 .lut_mask = 16'hEEFF;
defparam \sr~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~30 (
	.dataa(virtual_state_sdr),
	.datab(sr_27),
	.datac(\sr~28_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~30_combout ),
	.cout());
defparam \sr~30 .lut_mask = 16'hFEFF;
defparam \sr~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[33]~31 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[33]~31_combout ),
	.cout());
defparam \sr[33]~31 .lut_mask = 16'hFF7F;
defparam \sr[33]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~32 (
	.dataa(sr_35),
	.datab(virtual_state_sdr),
	.datac(monitor_error),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~32_combout ),
	.cout());
defparam \sr~32 .lut_mask = 16'hFFB8;
defparam \sr~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~33 (
	.dataa(break_readreg_27),
	.datab(MonDReg_27),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~33_combout ),
	.cout());
defparam \sr~33 .lut_mask = 16'hAACC;
defparam \sr~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~34 (
	.dataa(virtual_state_sdr),
	.datab(sr_29),
	.datac(\sr~33_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~34_combout ),
	.cout());
defparam \sr~34 .lut_mask = 16'hFEFF;
defparam \sr~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~35 (
	.dataa(break_readreg_26),
	.datab(MonDReg_26),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~35_combout ),
	.cout());
defparam \sr~35 .lut_mask = 16'hAACC;
defparam \sr~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~36 (
	.dataa(virtual_state_sdr),
	.datab(sr_28),
	.datac(\sr~35_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~36_combout ),
	.cout());
defparam \sr~36 .lut_mask = 16'hFEFF;
defparam \sr~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~37 (
	.dataa(break_readreg_24),
	.datab(MonDReg_24),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~37_combout ),
	.cout());
defparam \sr~37 .lut_mask = 16'hAACC;
defparam \sr~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~38 (
	.dataa(virtual_state_sdr),
	.datab(sr_26),
	.datac(\sr~37_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~38_combout ),
	.cout());
defparam \sr~38 .lut_mask = 16'hFEFF;
defparam \sr~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~39 (
	.dataa(break_readreg_16),
	.datab(MonDReg_16),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~39_combout ),
	.cout());
defparam \sr~39 .lut_mask = 16'hAACC;
defparam \sr~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~40 (
	.dataa(virtual_state_sdr),
	.datab(sr_18),
	.datac(\sr~39_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~40_combout ),
	.cout());
defparam \sr~40 .lut_mask = 16'hFEFF;
defparam \sr~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~41 (
	.dataa(break_readreg_20),
	.datab(MonDReg_20),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~41_combout ),
	.cout());
defparam \sr~41 .lut_mask = 16'hAACC;
defparam \sr~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~42 (
	.dataa(virtual_state_sdr),
	.datab(sr_22),
	.datac(\sr~41_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~42_combout ),
	.cout());
defparam \sr~42 .lut_mask = 16'hFEFF;
defparam \sr~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~43 (
	.dataa(break_readreg_19),
	.datab(MonDReg_19),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~43_combout ),
	.cout());
defparam \sr~43 .lut_mask = 16'hAACC;
defparam \sr~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~44 (
	.dataa(virtual_state_sdr),
	.datab(sr_21),
	.datac(\sr~43_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~44_combout ),
	.cout());
defparam \sr~44 .lut_mask = 16'hFEFF;
defparam \sr~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~45 (
	.dataa(break_readreg_5),
	.datab(MonDReg_5),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~45_combout ),
	.cout());
defparam \sr~45 .lut_mask = 16'hAACC;
defparam \sr~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~46 (
	.dataa(sr_7),
	.datab(virtual_state_sdr),
	.datac(\sr~45_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~46_combout ),
	.cout());
defparam \sr~46 .lut_mask = 16'hB8FF;
defparam \sr~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~47 (
	.dataa(break_readreg_28),
	.datab(MonDReg_28),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~47_combout ),
	.cout());
defparam \sr~47 .lut_mask = 16'hAACC;
defparam \sr~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~48 (
	.dataa(virtual_state_sdr),
	.datab(sr_30),
	.datac(\sr~47_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~48_combout ),
	.cout());
defparam \sr~48 .lut_mask = 16'hFEFF;
defparam \sr~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~49 (
	.dataa(break_readreg_29),
	.datab(MonDReg_29),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~49_combout ),
	.cout());
defparam \sr~49 .lut_mask = 16'hAACC;
defparam \sr~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~50 (
	.dataa(virtual_state_sdr),
	.datab(sr_31),
	.datac(\sr~49_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~50_combout ),
	.cout());
defparam \sr~50 .lut_mask = 16'hFEFF;
defparam \sr~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~52 (
	.dataa(break_readreg_31),
	.datab(MonDReg_31),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~52_combout ),
	.cout());
defparam \sr~52 .lut_mask = 16'hAACC;
defparam \sr~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~53 (
	.dataa(virtual_state_sdr),
	.datab(sr_33),
	.datac(\sr~52_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~53_combout ),
	.cout());
defparam \sr~53 .lut_mask = 16'hFEFF;
defparam \sr~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~54 (
	.dataa(sr_34),
	.datab(virtual_state_sdr),
	.datac(resetlatch),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~54_combout ),
	.cout());
defparam \sr~54 .lut_mask = 16'hFFB8;
defparam \sr~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~55 (
	.dataa(break_readreg_17),
	.datab(MonDReg_17),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~55_combout ),
	.cout());
defparam \sr~55 .lut_mask = 16'hAACC;
defparam \sr~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~56 (
	.dataa(virtual_state_sdr),
	.datab(sr_19),
	.datac(\sr~55_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~56_combout ),
	.cout());
defparam \sr~56 .lut_mask = 16'hFEFF;
defparam \sr~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~57 (
	.dataa(break_readreg_18),
	.datab(MonDReg_18),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~57_combout ),
	.cout());
defparam \sr~57 .lut_mask = 16'hAACC;
defparam \sr~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~58 (
	.dataa(virtual_state_sdr),
	.datab(sr_20),
	.datac(\sr~57_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~58_combout ),
	.cout());
defparam \sr~58 .lut_mask = 16'hFEFF;
defparam \sr~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~59 (
	.dataa(break_readreg_21),
	.datab(MonDReg_21),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~59_combout ),
	.cout());
defparam \sr~59 .lut_mask = 16'hAACC;
defparam \sr~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~60 (
	.dataa(virtual_state_sdr),
	.datab(sr_23),
	.datac(\sr~59_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~60_combout ),
	.cout());
defparam \sr~60 .lut_mask = 16'hFEFF;
defparam \sr~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~61 (
	.dataa(break_readreg_22),
	.datab(MonDReg_22),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~61_combout ),
	.cout());
defparam \sr~61 .lut_mask = 16'hAACC;
defparam \sr~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~62 (
	.dataa(virtual_state_sdr),
	.datab(sr_24),
	.datac(\sr~61_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~62_combout ),
	.cout());
defparam \sr~62 .lut_mask = 16'hFEFF;
defparam \sr~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~63 (
	.dataa(break_readreg_7),
	.datab(MonDReg_7),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~63_combout ),
	.cout());
defparam \sr~63 .lut_mask = 16'hAACC;
defparam \sr~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~64 (
	.dataa(sr_9),
	.datab(virtual_state_sdr),
	.datac(\sr~63_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~64_combout ),
	.cout());
defparam \sr~64 .lut_mask = 16'hB8FF;
defparam \sr~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~65 (
	.dataa(break_readreg_23),
	.datab(MonDReg_23),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~65_combout ),
	.cout());
defparam \sr~65 .lut_mask = 16'hAACC;
defparam \sr~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~66 (
	.dataa(virtual_state_sdr),
	.datab(sr_25),
	.datac(\sr~65_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~66_combout ),
	.cout());
defparam \sr~66 .lut_mask = 16'hFEFF;
defparam \sr~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~67 (
	.dataa(break_readreg_15),
	.datab(MonDReg_15),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~67_combout ),
	.cout());
defparam \sr~67 .lut_mask = 16'hAACC;
defparam \sr~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~68 (
	.dataa(virtual_state_sdr),
	.datab(sr_17),
	.datac(\sr~67_combout ),
	.datad(\sr~29_combout ),
	.cin(gnd),
	.combout(\sr~68_combout ),
	.cout());
defparam \sr~68 .lut_mask = 16'hFEFF;
defparam \sr~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~69 (
	.dataa(break_readreg_8),
	.datab(MonDReg_8),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~69_combout ),
	.cout());
defparam \sr~69 .lut_mask = 16'hAACC;
defparam \sr~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~70 (
	.dataa(sr_10),
	.datab(virtual_state_sdr),
	.datac(\sr~69_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~70_combout ),
	.cout());
defparam \sr~70 .lut_mask = 16'hB8FF;
defparam \sr~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~71 (
	.dataa(break_readreg_13),
	.datab(MonDReg_13),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~71_combout ),
	.cout());
defparam \sr~71 .lut_mask = 16'hAACC;
defparam \sr~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~72 (
	.dataa(sr_15),
	.datab(virtual_state_sdr),
	.datac(\sr~71_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~72_combout ),
	.cout());
defparam \sr~72 .lut_mask = 16'hB8FF;
defparam \sr~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~75 (
	.dataa(break_readreg_12),
	.datab(MonDReg_12),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~75_combout ),
	.cout());
defparam \sr~75 .lut_mask = 16'hAACC;
defparam \sr~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~76 (
	.dataa(sr_14),
	.datab(virtual_state_sdr),
	.datac(\sr~75_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~76_combout ),
	.cout());
defparam \sr~76 .lut_mask = 16'hB8FF;
defparam \sr~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~77 (
	.dataa(break_readreg_11),
	.datab(MonDReg_11),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~77_combout ),
	.cout());
defparam \sr~77 .lut_mask = 16'hAACC;
defparam \sr~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~78 (
	.dataa(sr_13),
	.datab(virtual_state_sdr),
	.datac(\sr~77_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~78_combout ),
	.cout());
defparam \sr~78 .lut_mask = 16'hB8FF;
defparam \sr~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~79 (
	.dataa(break_readreg_10),
	.datab(MonDReg_10),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~79_combout ),
	.cout());
defparam \sr~79 .lut_mask = 16'hAACC;
defparam \sr~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~80 (
	.dataa(sr_12),
	.datab(virtual_state_sdr),
	.datac(\sr~79_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~80_combout ),
	.cout());
defparam \sr~80 .lut_mask = 16'hB8FF;
defparam \sr~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~81 (
	.dataa(break_readreg_9),
	.datab(MonDReg_9),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~81_combout ),
	.cout());
defparam \sr~81 .lut_mask = 16'hAACC;
defparam \sr~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~82 (
	.dataa(sr_11),
	.datab(virtual_state_sdr),
	.datac(\sr~81_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~82_combout ),
	.cout());
defparam \sr~82 .lut_mask = 16'hB8FF;
defparam \sr~82 .sum_lutc_input = "datac";

endmodule

module niosII_altera_std_synchronizer_4 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_5 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_sld_virtual_jtag_basic_1 (
	virtual_state_cdr1,
	virtual_state_sdr,
	virtual_state_uir,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_cdr1;
output 	virtual_state_sdr;
output 	virtual_state_uir;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb virtual_state_cdr(
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(state_3),
	.datad(splitter_nodes_receive_1_3),
	.cin(gnd),
	.combout(virtual_state_cdr1),
	.cout());
defparam virtual_state_cdr.lut_mask = 16'hAFFF;
defparam virtual_state_cdr.sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_sdr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_sdr),
	.cout());
defparam \virtual_state_sdr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_sdr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_uir~0 (
	.dataa(virtual_ir_scan_reg),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_8),
	.datad(gnd),
	.cin(gnd),
	.combout(virtual_state_uir),
	.cout());
defparam \virtual_state_uir~0 .lut_mask = 16'hFEFE;
defparam \virtual_state_uir~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_udr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_8),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_udr),
	.cout());
defparam \virtual_state_udr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_udr~0 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_cpu_cpu_nios2_avalon_reg (
	wire_pll7_clk_0,
	r_sync_rst,
	address_8,
	ociram_wr_en,
	writedata_0,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	Equal0,
	Equal01,
	take_action_ocireg,
	oci_ienable_4,
	oci_ienable_3,
	oci_ienable_2,
	oci_ienable_1,
	oci_ienable_0,
	oci_single_step_mode1,
	writedata_1,
	writedata_4,
	writedata_3,
	writedata_2,
	Equal02,
	oci_reg_readdata,
	oci_ienable_23)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	address_8;
input 	ociram_wr_en;
input 	writedata_0;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
output 	Equal0;
output 	Equal01;
output 	take_action_ocireg;
output 	oci_ienable_4;
output 	oci_ienable_3;
output 	oci_ienable_2;
output 	oci_ienable_1;
output 	oci_ienable_0;
output 	oci_single_step_mode1;
input 	writedata_1;
input 	writedata_4;
input 	writedata_3;
input 	writedata_2;
output 	Equal02;
output 	oci_reg_readdata;
output 	oci_ienable_23;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \oci_ienable[4]~0_combout ;
wire \take_action_oci_intr_mask_reg~0_combout ;
wire \oci_ienable[3]~1_combout ;
wire \oci_ienable[2]~2_combout ;
wire \oci_ienable[1]~3_combout ;
wire \oci_ienable[0]~4_combout ;
wire \oci_single_step_mode~0_combout ;


cycloneive_lcell_comb \Equal0~0 (
	.dataa(address_8),
	.datab(address_5),
	.datac(address_6),
	.datad(address_7),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hBFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(address_1),
	.datab(address_2),
	.datac(address_3),
	.datad(address_4),
	.cin(gnd),
	.combout(Equal01),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_ocireg~0 (
	.dataa(ociram_wr_en),
	.datab(Equal0),
	.datac(Equal01),
	.datad(address_0),
	.cin(gnd),
	.combout(take_action_ocireg),
	.cout());
defparam \take_action_ocireg~0 .lut_mask = 16'hFEFF;
defparam \take_action_ocireg~0 .sum_lutc_input = "datac";

dffeas \oci_ienable[4] (
	.clk(wire_pll7_clk_0),
	.d(\oci_ienable[4]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_4),
	.prn(vcc));
defparam \oci_ienable[4] .is_wysiwyg = "true";
defparam \oci_ienable[4] .power_up = "low";

dffeas \oci_ienable[3] (
	.clk(wire_pll7_clk_0),
	.d(\oci_ienable[3]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_3),
	.prn(vcc));
defparam \oci_ienable[3] .is_wysiwyg = "true";
defparam \oci_ienable[3] .power_up = "low";

dffeas \oci_ienable[2] (
	.clk(wire_pll7_clk_0),
	.d(\oci_ienable[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_2),
	.prn(vcc));
defparam \oci_ienable[2] .is_wysiwyg = "true";
defparam \oci_ienable[2] .power_up = "low";

dffeas \oci_ienable[1] (
	.clk(wire_pll7_clk_0),
	.d(\oci_ienable[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_1),
	.prn(vcc));
defparam \oci_ienable[1] .is_wysiwyg = "true";
defparam \oci_ienable[1] .power_up = "low";

dffeas \oci_ienable[0] (
	.clk(wire_pll7_clk_0),
	.d(\oci_ienable[0]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_0),
	.prn(vcc));
defparam \oci_ienable[0] .is_wysiwyg = "true";
defparam \oci_ienable[0] .power_up = "low";

dffeas oci_single_step_mode(
	.clk(wire_pll7_clk_0),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(Equal0),
	.datab(Equal01),
	.datac(gnd),
	.datad(address_0),
	.cin(gnd),
	.combout(Equal02),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_reg_readdata~0 (
	.dataa(address_0),
	.datab(Equal0),
	.datac(Equal01),
	.datad(oci_ienable_4),
	.cin(gnd),
	.combout(oci_reg_readdata),
	.cout());
defparam \oci_reg_readdata~0 .lut_mask = 16'hFEFF;
defparam \oci_reg_readdata~0 .sum_lutc_input = "datac";

dffeas \oci_ienable[23] (
	.clk(wire_pll7_clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_23),
	.prn(vcc));
defparam \oci_ienable[23] .is_wysiwyg = "true";
defparam \oci_ienable[23] .power_up = "low";

cycloneive_lcell_comb \oci_ienable[4]~0 (
	.dataa(writedata_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[4]~0_combout ),
	.cout());
defparam \oci_ienable[4]~0 .lut_mask = 16'h5555;
defparam \oci_ienable[4]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_oci_intr_mask_reg~0 (
	.dataa(ociram_wr_en),
	.datab(address_0),
	.datac(Equal0),
	.datad(Equal01),
	.cin(gnd),
	.combout(\take_action_oci_intr_mask_reg~0_combout ),
	.cout());
defparam \take_action_oci_intr_mask_reg~0 .lut_mask = 16'hFFFE;
defparam \take_action_oci_intr_mask_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_ienable[3]~1 (
	.dataa(writedata_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[3]~1_combout ),
	.cout());
defparam \oci_ienable[3]~1 .lut_mask = 16'h5555;
defparam \oci_ienable[3]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_ienable[2]~2 (
	.dataa(writedata_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[2]~2_combout ),
	.cout());
defparam \oci_ienable[2]~2 .lut_mask = 16'h5555;
defparam \oci_ienable[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_ienable[1]~3 (
	.dataa(writedata_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[1]~3_combout ),
	.cout());
defparam \oci_ienable[1]~3 .lut_mask = 16'h5555;
defparam \oci_ienable[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_ienable[0]~4 (
	.dataa(writedata_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[0]~4_combout ),
	.cout());
defparam \oci_ienable[0]~4 .lut_mask = 16'h5555;
defparam \oci_ienable[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_single_step_mode~0 (
	.dataa(writedata_3),
	.datab(oci_single_step_mode1),
	.datac(gnd),
	.datad(take_action_ocireg),
	.cin(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.cout());
defparam \oci_single_step_mode~0 .lut_mask = 16'hAACC;
defparam \oci_single_step_mode~0 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_cpu_cpu_nios2_oci_break (
	wire_pll7_clk_0,
	break_readreg_0,
	break_readreg_1,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_0,
	ir_1,
	enable_action_strobe,
	jdo_3,
	break_readreg_2,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_17,
	jdo_21,
	jdo_20,
	break_readreg_3,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_19,
	jdo_18,
	break_readreg_4,
	jdo_6,
	break_readreg_25,
	break_readreg_27,
	break_readreg_26,
	break_readreg_24,
	break_readreg_16,
	break_readreg_20,
	break_readreg_19,
	jdo_23,
	break_readreg_5,
	jdo_7,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	jdo_24,
	break_readreg_17,
	jdo_16,
	jdo_22,
	break_readreg_18,
	break_readreg_21,
	break_readreg_6,
	jdo_8,
	jdo_14,
	jdo_15,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_22,
	break_readreg_7,
	break_readreg_23,
	break_readreg_15,
	break_readreg_8,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	break_readreg_0;
output 	break_readreg_1;
input 	jdo_0;
input 	jdo_36;
input 	jdo_37;
input 	ir_0;
input 	ir_1;
input 	enable_action_strobe;
input 	jdo_3;
output 	break_readreg_2;
input 	jdo_1;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	jdo_25;
input 	jdo_17;
input 	jdo_21;
input 	jdo_20;
output 	break_readreg_3;
input 	jdo_2;
input 	jdo_5;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_19;
input 	jdo_18;
output 	break_readreg_4;
input 	jdo_6;
output 	break_readreg_25;
output 	break_readreg_27;
output 	break_readreg_26;
output 	break_readreg_24;
output 	break_readreg_16;
output 	break_readreg_20;
output 	break_readreg_19;
input 	jdo_23;
output 	break_readreg_5;
input 	jdo_7;
output 	break_readreg_28;
output 	break_readreg_29;
output 	break_readreg_30;
output 	break_readreg_31;
input 	jdo_24;
output 	break_readreg_17;
input 	jdo_16;
input 	jdo_22;
output 	break_readreg_18;
output 	break_readreg_21;
output 	break_readreg_6;
input 	jdo_8;
input 	jdo_14;
input 	jdo_15;
input 	jdo_13;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;
output 	break_readreg_22;
output 	break_readreg_7;
output 	break_readreg_23;
output 	break_readreg_15;
output 	break_readreg_8;
output 	break_readreg_13;
output 	break_readreg_14;
output 	break_readreg_12;
output 	break_readreg_11;
output 	break_readreg_10;
output 	break_readreg_9;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg~0_combout ;
wire \break_readreg[31]~1_combout ;
wire \break_readreg~2_combout ;
wire \break_readreg~3_combout ;
wire \break_readreg~4_combout ;
wire \break_readreg~5_combout ;
wire \break_readreg~6_combout ;
wire \break_readreg~7_combout ;
wire \break_readreg~8_combout ;
wire \break_readreg~9_combout ;
wire \break_readreg~10_combout ;
wire \break_readreg~11_combout ;
wire \break_readreg~12_combout ;
wire \break_readreg~13_combout ;
wire \break_readreg~14_combout ;
wire \break_readreg~15_combout ;
wire \break_readreg~16_combout ;
wire \break_readreg~17_combout ;
wire \break_readreg~18_combout ;
wire \break_readreg~19_combout ;
wire \break_readreg~20_combout ;
wire \break_readreg~21_combout ;
wire \break_readreg~22_combout ;
wire \break_readreg~23_combout ;
wire \break_readreg~24_combout ;
wire \break_readreg~25_combout ;
wire \break_readreg~26_combout ;
wire \break_readreg~27_combout ;
wire \break_readreg~28_combout ;
wire \break_readreg~29_combout ;
wire \break_readreg~30_combout ;
wire \break_readreg~31_combout ;
wire \break_readreg~32_combout ;


dffeas \break_readreg[0] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(wire_pll7_clk_0),
	.d(\break_readreg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[31]~1_combout ),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

cycloneive_lcell_comb \break_readreg~0 (
	.dataa(jdo_0),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(gnd),
	.cin(gnd),
	.combout(\break_readreg~0_combout ),
	.cout());
defparam \break_readreg~0 .lut_mask = 16'hFEFE;
defparam \break_readreg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg[31]~1 (
	.dataa(ir_0),
	.datab(gnd),
	.datac(ir_1),
	.datad(enable_action_strobe),
	.cin(gnd),
	.combout(\break_readreg[31]~1_combout ),
	.cout());
defparam \break_readreg[31]~1 .lut_mask = 16'hFFF5;
defparam \break_readreg[31]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~2 (
	.dataa(jdo_1),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(gnd),
	.cin(gnd),
	.combout(\break_readreg~2_combout ),
	.cout());
defparam \break_readreg~2 .lut_mask = 16'hFEFE;
defparam \break_readreg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~3 (
	.dataa(jdo_2),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(gnd),
	.cin(gnd),
	.combout(\break_readreg~3_combout ),
	.cout());
defparam \break_readreg~3 .lut_mask = 16'hFEFE;
defparam \break_readreg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~4 (
	.dataa(jdo_3),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~4_combout ),
	.cout());
defparam \break_readreg~4 .lut_mask = 16'hFEFF;
defparam \break_readreg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~5 (
	.dataa(jdo_4),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~5_combout ),
	.cout());
defparam \break_readreg~5 .lut_mask = 16'hFEFF;
defparam \break_readreg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~6 (
	.dataa(jdo_25),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~6_combout ),
	.cout());
defparam \break_readreg~6 .lut_mask = 16'hFEFF;
defparam \break_readreg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~7 (
	.dataa(jdo_27),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~7_combout ),
	.cout());
defparam \break_readreg~7 .lut_mask = 16'hFEFF;
defparam \break_readreg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~8 (
	.dataa(jdo_26),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~8_combout ),
	.cout());
defparam \break_readreg~8 .lut_mask = 16'hFEFF;
defparam \break_readreg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~9 (
	.dataa(jdo_24),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~9_combout ),
	.cout());
defparam \break_readreg~9 .lut_mask = 16'hFEFF;
defparam \break_readreg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~10 (
	.dataa(jdo_16),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~10_combout ),
	.cout());
defparam \break_readreg~10 .lut_mask = 16'hFEFF;
defparam \break_readreg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~11 (
	.dataa(jdo_20),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~11_combout ),
	.cout());
defparam \break_readreg~11 .lut_mask = 16'hFEFF;
defparam \break_readreg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~12 (
	.dataa(jdo_19),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~12_combout ),
	.cout());
defparam \break_readreg~12 .lut_mask = 16'hFEFF;
defparam \break_readreg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~13 (
	.dataa(jdo_5),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~13_combout ),
	.cout());
defparam \break_readreg~13 .lut_mask = 16'hFEFF;
defparam \break_readreg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~14 (
	.dataa(jdo_28),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~14_combout ),
	.cout());
defparam \break_readreg~14 .lut_mask = 16'hFEFF;
defparam \break_readreg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~15 (
	.dataa(jdo_29),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~15_combout ),
	.cout());
defparam \break_readreg~15 .lut_mask = 16'hFEFF;
defparam \break_readreg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~16 (
	.dataa(jdo_30),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~16_combout ),
	.cout());
defparam \break_readreg~16 .lut_mask = 16'hFEFF;
defparam \break_readreg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~17 (
	.dataa(jdo_31),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~17_combout ),
	.cout());
defparam \break_readreg~17 .lut_mask = 16'hFEFF;
defparam \break_readreg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~18 (
	.dataa(jdo_17),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~18_combout ),
	.cout());
defparam \break_readreg~18 .lut_mask = 16'hFEFF;
defparam \break_readreg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~19 (
	.dataa(jdo_18),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~19_combout ),
	.cout());
defparam \break_readreg~19 .lut_mask = 16'hFEFF;
defparam \break_readreg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~20 (
	.dataa(jdo_21),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~20_combout ),
	.cout());
defparam \break_readreg~20 .lut_mask = 16'hFEFF;
defparam \break_readreg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~21 (
	.dataa(jdo_6),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~21_combout ),
	.cout());
defparam \break_readreg~21 .lut_mask = 16'hFEFF;
defparam \break_readreg~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~22 (
	.dataa(jdo_22),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~22_combout ),
	.cout());
defparam \break_readreg~22 .lut_mask = 16'hFEFF;
defparam \break_readreg~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~23 (
	.dataa(jdo_7),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~23_combout ),
	.cout());
defparam \break_readreg~23 .lut_mask = 16'hFEFF;
defparam \break_readreg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~24 (
	.dataa(jdo_23),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~24_combout ),
	.cout());
defparam \break_readreg~24 .lut_mask = 16'hFEFF;
defparam \break_readreg~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~25 (
	.dataa(jdo_15),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~25_combout ),
	.cout());
defparam \break_readreg~25 .lut_mask = 16'hFEFF;
defparam \break_readreg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~26 (
	.dataa(jdo_8),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~26_combout ),
	.cout());
defparam \break_readreg~26 .lut_mask = 16'hFEFF;
defparam \break_readreg~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~27 (
	.dataa(jdo_13),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~27_combout ),
	.cout());
defparam \break_readreg~27 .lut_mask = 16'hFEFF;
defparam \break_readreg~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~28 (
	.dataa(jdo_14),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~28_combout ),
	.cout());
defparam \break_readreg~28 .lut_mask = 16'hFEFF;
defparam \break_readreg~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~29 (
	.dataa(jdo_12),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~29_combout ),
	.cout());
defparam \break_readreg~29 .lut_mask = 16'hFEFF;
defparam \break_readreg~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~30 (
	.dataa(jdo_11),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~30_combout ),
	.cout());
defparam \break_readreg~30 .lut_mask = 16'hFEFF;
defparam \break_readreg~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~31 (
	.dataa(jdo_10),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~31_combout ),
	.cout());
defparam \break_readreg~31 .lut_mask = 16'hFEFF;
defparam \break_readreg~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~32 (
	.dataa(jdo_9),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[31]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~32_combout ),
	.cout());
defparam \break_readreg~32 .lut_mask = 16'hFEFF;
defparam \break_readreg~32 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_cpu_cpu_nios2_oci_debug (
	wire_pll7_clk_0,
	jtag_break1,
	r_sync_rst,
	take_action_ocimem_a,
	monitor_ready1,
	jdo_34,
	writedata_0,
	take_action_ocireg,
	jdo_25,
	jdo_21,
	jdo_20,
	take_action_ocimem_a1,
	writedata_1,
	jdo_19,
	jdo_18,
	monitor_error1,
	monitor_go1,
	resetrequest1,
	jdo_23,
	resetlatch1,
	jdo_24,
	jdo_22,
	state_1)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	jtag_break1;
input 	r_sync_rst;
input 	take_action_ocimem_a;
output 	monitor_ready1;
input 	jdo_34;
input 	writedata_0;
input 	take_action_ocireg;
input 	jdo_25;
input 	jdo_21;
input 	jdo_20;
input 	take_action_ocimem_a1;
input 	writedata_1;
input 	jdo_19;
input 	jdo_18;
output 	monitor_error1;
output 	monitor_go1;
output 	resetrequest1;
input 	jdo_23;
output 	resetlatch1;
input 	jdo_24;
input 	jdo_22;
input 	state_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \jtag_break~1_combout ;
wire \always1~0_combout ;
wire \monitor_ready~0_combout ;
wire \monitor_error~0_combout ;
wire \monitor_go~0_combout ;
wire \resetlatch~0_combout ;


niosII_altera_std_synchronizer_6 the_altera_std_synchronizer(
	.clk(wire_pll7_clk_0),
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ));

dffeas jtag_break(
	.clk(wire_pll7_clk_0),
	.d(\jtag_break~0_combout ),
	.asdata(\jtag_break~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_ready(
	.clk(wire_pll7_clk_0),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas monitor_error(
	.clk(wire_pll7_clk_0),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas monitor_go(
	.clk(wire_pll7_clk_0),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

dffeas resetrequest(
	.clk(wire_pll7_clk_0),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(resetrequest1),
	.prn(vcc));
defparam resetrequest.is_wysiwyg = "true";
defparam resetrequest.power_up = "low";

dffeas resetlatch(
	.clk(wire_pll7_clk_0),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

cycloneive_lcell_comb \break_on_reset~0 (
	.dataa(jdo_19),
	.datab(\break_on_reset~q ),
	.datac(gnd),
	.datad(jdo_18),
	.cin(gnd),
	.combout(\break_on_reset~0_combout ),
	.cout());
defparam \break_on_reset~0 .lut_mask = 16'hEEFF;
defparam \break_on_reset~0 .sum_lutc_input = "datac";

dffeas break_on_reset(
	.clk(wire_pll7_clk_0),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cycloneive_lcell_comb \jtag_break~0 (
	.dataa(jtag_break1),
	.datab(\break_on_reset~q ),
	.datac(gnd),
	.datad(\the_altera_std_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\jtag_break~0_combout ),
	.cout());
defparam \jtag_break~0 .lut_mask = 16'hAACC;
defparam \jtag_break~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_break~1 (
	.dataa(jdo_21),
	.datab(jtag_break1),
	.datac(gnd),
	.datad(jdo_20),
	.cin(gnd),
	.combout(\jtag_break~1_combout ),
	.cout());
defparam \jtag_break~1 .lut_mask = 16'hEEFF;
defparam \jtag_break~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(take_action_ocimem_a),
	.datab(jdo_34),
	.datac(jdo_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hFDFD;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_ready~0 (
	.dataa(monitor_ready1),
	.datab(writedata_0),
	.datac(take_action_ocireg),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_ready~0_combout ),
	.cout());
defparam \monitor_ready~0 .lut_mask = 16'hFEFF;
defparam \monitor_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_error~0 (
	.dataa(monitor_error1),
	.datab(take_action_ocireg),
	.datac(writedata_1),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_error~0_combout ),
	.cout());
defparam \monitor_error~0 .lut_mask = 16'hFEFF;
defparam \monitor_error~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_go~0 (
	.dataa(take_action_ocimem_a1),
	.datab(jdo_23),
	.datac(monitor_go1),
	.datad(state_1),
	.cin(gnd),
	.combout(\monitor_go~0_combout ),
	.cout());
defparam \monitor_go~0 .lut_mask = 16'hFEFF;
defparam \monitor_go~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \resetlatch~0 (
	.dataa(resetlatch1),
	.datab(\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(jdo_24),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\resetlatch~0_combout ),
	.cout());
defparam \resetlatch~0 .lut_mask = 16'hEFFF;
defparam \resetlatch~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_std_synchronizer_6 (
	clk,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_niosII_cpu_cpu_nios2_ocimem (
	wire_pll7_clk_0,
	MonDReg_0,
	MonDReg_1,
	q_a_0,
	q_a_1,
	MonDReg_3,
	q_a_2,
	q_a_3,
	q_a_4,
	MonDReg_4,
	MonDReg_25,
	MonDReg_26,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_21,
	q_a_30,
	q_a_29,
	q_a_28,
	q_a_27,
	q_a_26,
	q_a_25,
	q_a_24,
	q_a_23,
	q_a_22,
	q_a_20,
	q_a_19,
	q_a_18,
	q_a_17,
	MonDReg_5,
	MonDReg_29,
	MonDReg_11,
	MonDReg_12,
	q_a_31,
	MonDReg_9,
	MonDReg_8,
	MonDReg_18,
	waitrequest1,
	jdo_3,
	take_action_ocimem_b,
	take_no_action_ocimem_a,
	write,
	address_8,
	read,
	MonDReg_2,
	jdo_4,
	jdo_26,
	jdo_34,
	take_action_ocimem_a,
	jdo_28,
	jdo_27,
	debugaccess,
	ociram_wr_en,
	r_early_rst,
	writedata_0,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	byteenable_0,
	jdo_25,
	jdo_17,
	jdo_21,
	jdo_20,
	jdo_5,
	writedata_1,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	writedata_4,
	writedata_3,
	writedata_2,
	jdo_19,
	jdo_18,
	jdo_6,
	MonDReg_27,
	MonDReg_24,
	MonDReg_16,
	MonDReg_20,
	MonDReg_19,
	jdo_23,
	jdo_7,
	MonDReg_28,
	MonDReg_30,
	MonDReg_31,
	jdo_24,
	MonDReg_17,
	jdo_16,
	writedata_11,
	byteenable_1,
	MonDReg_13,
	writedata_13,
	writedata_16,
	byteenable_2,
	writedata_12,
	writedata_5,
	MonDReg_14,
	writedata_14,
	MonDReg_15,
	writedata_15,
	MonDReg_10,
	writedata_10,
	writedata_9,
	writedata_8,
	MonDReg_7,
	writedata_7,
	MonDReg_6,
	writedata_6,
	MonDReg_21,
	writedata_21,
	writedata_30,
	byteenable_3,
	writedata_29,
	writedata_28,
	writedata_27,
	writedata_26,
	writedata_25,
	writedata_24,
	MonDReg_23,
	writedata_23,
	MonDReg_22,
	writedata_22,
	writedata_20,
	writedata_19,
	writedata_18,
	writedata_17,
	jdo_22,
	jdo_8,
	jdo_14,
	jdo_15,
	jdo_13,
	writedata_31,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	MonDReg_0;
output 	MonDReg_1;
output 	q_a_0;
output 	q_a_1;
output 	MonDReg_3;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	MonDReg_4;
output 	MonDReg_25;
output 	MonDReg_26;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_10;
output 	q_a_9;
output 	q_a_8;
output 	q_a_7;
output 	q_a_6;
output 	q_a_21;
output 	q_a_30;
output 	q_a_29;
output 	q_a_28;
output 	q_a_27;
output 	q_a_26;
output 	q_a_25;
output 	q_a_24;
output 	q_a_23;
output 	q_a_22;
output 	q_a_20;
output 	q_a_19;
output 	q_a_18;
output 	q_a_17;
output 	MonDReg_5;
output 	MonDReg_29;
output 	MonDReg_11;
output 	MonDReg_12;
output 	q_a_31;
output 	MonDReg_9;
output 	MonDReg_8;
output 	MonDReg_18;
output 	waitrequest1;
input 	jdo_3;
input 	take_action_ocimem_b;
input 	take_no_action_ocimem_a;
input 	write;
input 	address_8;
input 	read;
output 	MonDReg_2;
input 	jdo_4;
input 	jdo_26;
input 	jdo_34;
input 	take_action_ocimem_a;
input 	jdo_28;
input 	jdo_27;
input 	debugaccess;
output 	ociram_wr_en;
input 	r_early_rst;
input 	writedata_0;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
input 	byteenable_0;
input 	jdo_25;
input 	jdo_17;
input 	jdo_21;
input 	jdo_20;
input 	jdo_5;
input 	writedata_1;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_32;
input 	jdo_33;
input 	writedata_4;
input 	writedata_3;
input 	writedata_2;
input 	jdo_19;
input 	jdo_18;
input 	jdo_6;
output 	MonDReg_27;
output 	MonDReg_24;
output 	MonDReg_16;
output 	MonDReg_20;
output 	MonDReg_19;
input 	jdo_23;
input 	jdo_7;
output 	MonDReg_28;
output 	MonDReg_30;
output 	MonDReg_31;
input 	jdo_24;
output 	MonDReg_17;
input 	jdo_16;
input 	writedata_11;
input 	byteenable_1;
output 	MonDReg_13;
input 	writedata_13;
input 	writedata_16;
input 	byteenable_2;
input 	writedata_12;
input 	writedata_5;
output 	MonDReg_14;
input 	writedata_14;
output 	MonDReg_15;
input 	writedata_15;
output 	MonDReg_10;
input 	writedata_10;
input 	writedata_9;
input 	writedata_8;
output 	MonDReg_7;
input 	writedata_7;
output 	MonDReg_6;
input 	writedata_6;
output 	MonDReg_21;
input 	writedata_21;
input 	writedata_30;
input 	byteenable_3;
input 	writedata_29;
input 	writedata_28;
input 	writedata_27;
input 	writedata_26;
input 	writedata_25;
input 	writedata_24;
output 	MonDReg_23;
input 	writedata_23;
output 	MonDReg_22;
input 	writedata_22;
input 	writedata_20;
input 	writedata_19;
input 	writedata_18;
input 	writedata_17;
input 	jdo_22;
input 	jdo_8;
input 	jdo_14;
input 	jdo_15;
input 	jdo_13;
input 	writedata_31;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_ram_wr~q ;
wire \ociram_wr_en~1_combout ;
wire \ociram_reset_req~combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[3]~3_combout ;
wire \ociram_wr_data[4]~4_combout ;
wire \ociram_wr_data[11]~5_combout ;
wire \ociram_byteenable[1]~1_combout ;
wire \ociram_wr_data[13]~6_combout ;
wire \ociram_wr_data[16]~7_combout ;
wire \ociram_byteenable[2]~2_combout ;
wire \ociram_wr_data[12]~8_combout ;
wire \ociram_wr_data[5]~9_combout ;
wire \ociram_wr_data[14]~10_combout ;
wire \ociram_wr_data[15]~11_combout ;
wire \ociram_wr_data[10]~12_combout ;
wire \ociram_wr_data[9]~13_combout ;
wire \ociram_wr_data[8]~14_combout ;
wire \ociram_wr_data[7]~15_combout ;
wire \ociram_wr_data[6]~16_combout ;
wire \ociram_wr_data[21]~17_combout ;
wire \ociram_wr_data[30]~18_combout ;
wire \ociram_byteenable[3]~3_combout ;
wire \ociram_wr_data[29]~19_combout ;
wire \ociram_wr_data[28]~20_combout ;
wire \ociram_wr_data[27]~21_combout ;
wire \ociram_wr_data[26]~22_combout ;
wire \ociram_wr_data[25]~23_combout ;
wire \ociram_wr_data[24]~24_combout ;
wire \ociram_wr_data[23]~25_combout ;
wire \ociram_wr_data[22]~26_combout ;
wire \ociram_wr_data[20]~27_combout ;
wire \ociram_wr_data[19]~28_combout ;
wire \ociram_wr_data[18]~29_combout ;
wire \ociram_wr_data[17]~30_combout ;
wire \ociram_wr_data[31]~31_combout ;
wire \MonARegAddrInc[0]~0_combout ;
wire \MonAReg~0_combout ;
wire \MonAReg[2]~q ;
wire \MonARegAddrInc[0]~1 ;
wire \MonARegAddrInc[1]~2_combout ;
wire \MonAReg~2_combout ;
wire \MonAReg[3]~q ;
wire \MonARegAddrInc[1]~3 ;
wire \MonARegAddrInc[2]~4_combout ;
wire \MonAReg~1_combout ;
wire \MonAReg[4]~q ;
wire \Equal0~0_combout ;
wire \jtag_ram_access~0_combout ;
wire \MonAReg[10]~q ;
wire \MonARegAddrInc[2]~5 ;
wire \MonARegAddrInc[3]~6_combout ;
wire \MonAReg~3_combout ;
wire \MonAReg[5]~q ;
wire \MonARegAddrInc[3]~7 ;
wire \MonARegAddrInc[4]~8_combout ;
wire \MonAReg~4_combout ;
wire \MonAReg[6]~q ;
wire \MonARegAddrInc[4]~9 ;
wire \MonARegAddrInc[5]~10_combout ;
wire \MonAReg~5_combout ;
wire \MonAReg[7]~q ;
wire \MonARegAddrInc[5]~11 ;
wire \MonARegAddrInc[6]~12_combout ;
wire \MonAReg~6_combout ;
wire \MonAReg[8]~q ;
wire \MonARegAddrInc[6]~13 ;
wire \MonARegAddrInc[7]~14_combout ;
wire \MonAReg~7_combout ;
wire \MonAReg[9]~q ;
wire \MonARegAddrInc[7]~15 ;
wire \MonARegAddrInc[8]~16_combout ;
wire \jtag_ram_rd~0_combout ;
wire \jtag_ram_rd~1_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[0]~0_combout ;
wire \jtag_rd~0_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~13_combout ;
wire \MonDReg[1]~1_combout ;
wire \MonDReg[3]~2_combout ;
wire \MonDReg[4]~3_combout ;
wire \Equal0~1_combout ;
wire \MonDReg[25]~5_combout ;
wire \Equal0~2_combout ;
wire \MonDReg[26]~4_combout ;
wire \MonDReg[5]~6_combout ;
wire \Equal0~3_combout ;
wire \MonDReg[29]~7_combout ;
wire \MonDReg[11]~8_combout ;
wire \Equal0~4_combout ;
wire \MonDReg[12]~9_combout ;
wire \MonDReg[9]~10_combout ;
wire \MonDReg~28_combout ;
wire \MonDReg[8]~11_combout ;
wire \Equal0~5_combout ;
wire \MonDReg[18]~12_combout ;
wire \jtag_ram_access~1_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~1_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~14_combout ;
wire \MonDReg~15_combout ;
wire \MonDReg~16_combout ;
wire \MonDReg~17_combout ;
wire \MonDReg~18_combout ;
wire \MonDReg~19_combout ;
wire \MonDReg~20_combout ;
wire \MonDReg~21_combout ;
wire \MonDReg~22_combout ;
wire \MonDReg~23_combout ;
wire \MonDReg~24_combout ;
wire \MonDReg~25_combout ;
wire \MonDReg~26_combout ;
wire \MonDReg~27_combout ;
wire \MonDReg~29_combout ;
wire \MonDReg~30_combout ;
wire \MonDReg~31_combout ;
wire \MonDReg~32_combout ;
wire \MonDReg~33_combout ;


niosII_niosII_cpu_cpu_ociram_sp_ram_module niosII_cpu_cpu_ociram_sp_ram(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_11(q_a_11),
	.q_a_13(q_a_13),
	.q_a_16(q_a_16),
	.q_a_12(q_a_12),
	.q_a_5(q_a_5),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_10(q_a_10),
	.q_a_9(q_a_9),
	.q_a_8(q_a_8),
	.q_a_7(q_a_7),
	.q_a_6(q_a_6),
	.q_a_21(q_a_21),
	.q_a_30(q_a_30),
	.q_a_29(q_a_29),
	.q_a_28(q_a_28),
	.q_a_27(q_a_27),
	.q_a_26(q_a_26),
	.q_a_25(q_a_25),
	.q_a_24(q_a_24),
	.q_a_23(q_a_23),
	.q_a_22(q_a_22),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.q_a_18(q_a_18),
	.q_a_17(q_a_17),
	.q_a_31(q_a_31),
	.ociram_wr_en(\ociram_wr_en~1_combout ),
	.ociram_reset_req(\ociram_reset_req~combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~3_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~4_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~5_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~1_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~6_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~7_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~2_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~8_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~9_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~10_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~11_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~12_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~13_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~14_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~15_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~16_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~17_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~18_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~3_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~19_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~20_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~21_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~22_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~23_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~24_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~25_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~26_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~27_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~28_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~29_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~30_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~31_combout ));

dffeas jtag_ram_wr(
	.clk(wire_pll7_clk_0),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_ocimem_a),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cycloneive_lcell_comb \ociram_wr_en~1 (
	.dataa(\jtag_ram_wr~q ),
	.datab(\jtag_ram_access~q ),
	.datac(ociram_wr_en),
	.datad(address_8),
	.cin(gnd),
	.combout(\ociram_wr_en~1_combout ),
	.cout());
defparam \ociram_wr_en~1 .lut_mask = 16'hB8FF;
defparam \ociram_wr_en~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb ociram_reset_req(
	.dataa(r_early_rst),
	.datab(gnd),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_reset_req~combout ),
	.cout());
defparam ociram_reset_req.lut_mask = 16'hFF55;
defparam ociram_reset_req.sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(MonDReg_0),
	.datab(writedata_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.cout());
defparam \ociram_wr_data[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(address_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.cout());
defparam \ociram_addr[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_addr[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[1]~1 (
	.dataa(\MonAReg[3]~q ),
	.datab(address_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.cout());
defparam \ociram_addr[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_addr[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[2]~2 (
	.dataa(\MonAReg[4]~q ),
	.datab(address_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.cout());
defparam \ociram_addr[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_addr[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[3]~3 (
	.dataa(\MonAReg[5]~q ),
	.datab(address_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.cout());
defparam \ociram_addr[3]~3 .lut_mask = 16'hAACC;
defparam \ociram_addr[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[4]~4 (
	.dataa(\MonAReg[6]~q ),
	.datab(address_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.cout());
defparam \ociram_addr[4]~4 .lut_mask = 16'hAACC;
defparam \ociram_addr[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[5]~5 (
	.dataa(\MonAReg[7]~q ),
	.datab(address_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.cout());
defparam \ociram_addr[5]~5 .lut_mask = 16'hAACC;
defparam \ociram_addr[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[6]~6 (
	.dataa(\MonAReg[8]~q ),
	.datab(address_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.cout());
defparam \ociram_addr[6]~6 .lut_mask = 16'hAACC;
defparam \ociram_addr[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[7]~7 (
	.dataa(\MonAReg[9]~q ),
	.datab(address_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.cout());
defparam \ociram_addr[7]~7 .lut_mask = 16'hAACC;
defparam \ociram_addr[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.cout());
defparam \ociram_byteenable[0]~0 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(MonDReg_1),
	.datab(writedata_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.cout());
defparam \ociram_wr_data[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_wr~0 (
	.dataa(\MonARegAddrInc[8]~16_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.cout());
defparam \jtag_ram_wr~0 .lut_mask = 16'hFF55;
defparam \jtag_ram_wr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(MonDReg_2),
	.datab(writedata_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.cout());
defparam \ociram_wr_data[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[3]~3 (
	.dataa(MonDReg_3),
	.datab(writedata_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[3]~3_combout ),
	.cout());
defparam \ociram_wr_data[3]~3 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[4]~4 (
	.dataa(MonDReg_4),
	.datab(writedata_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[4]~4_combout ),
	.cout());
defparam \ociram_wr_data[4]~4 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[11]~5 (
	.dataa(MonDReg_11),
	.datab(writedata_11),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[11]~5_combout ),
	.cout());
defparam \ociram_wr_data[11]~5 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[11]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[1]~1 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[1]~1_combout ),
	.cout());
defparam \ociram_byteenable[1]~1 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[13]~6 (
	.dataa(MonDReg_13),
	.datab(writedata_13),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[13]~6_combout ),
	.cout());
defparam \ociram_wr_data[13]~6 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[13]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[16]~7 (
	.dataa(MonDReg_16),
	.datab(writedata_16),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[16]~7_combout ),
	.cout());
defparam \ociram_wr_data[16]~7 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[16]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[2]~2 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[2]~2_combout ),
	.cout());
defparam \ociram_byteenable[2]~2 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[12]~8 (
	.dataa(MonDReg_12),
	.datab(writedata_12),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[12]~8_combout ),
	.cout());
defparam \ociram_wr_data[12]~8 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[12]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[5]~9 (
	.dataa(MonDReg_5),
	.datab(writedata_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[5]~9_combout ),
	.cout());
defparam \ociram_wr_data[5]~9 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[5]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[14]~10 (
	.dataa(MonDReg_14),
	.datab(writedata_14),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[14]~10_combout ),
	.cout());
defparam \ociram_wr_data[14]~10 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[14]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[15]~11 (
	.dataa(MonDReg_15),
	.datab(writedata_15),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[15]~11_combout ),
	.cout());
defparam \ociram_wr_data[15]~11 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[15]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[10]~12 (
	.dataa(MonDReg_10),
	.datab(writedata_10),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[10]~12_combout ),
	.cout());
defparam \ociram_wr_data[10]~12 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[10]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[9]~13 (
	.dataa(MonDReg_9),
	.datab(writedata_9),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[9]~13_combout ),
	.cout());
defparam \ociram_wr_data[9]~13 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[9]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[8]~14 (
	.dataa(MonDReg_8),
	.datab(writedata_8),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[8]~14_combout ),
	.cout());
defparam \ociram_wr_data[8]~14 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[8]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[7]~15 (
	.dataa(MonDReg_7),
	.datab(writedata_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[7]~15_combout ),
	.cout());
defparam \ociram_wr_data[7]~15 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[7]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[6]~16 (
	.dataa(MonDReg_6),
	.datab(writedata_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[6]~16_combout ),
	.cout());
defparam \ociram_wr_data[6]~16 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[6]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[21]~17 (
	.dataa(MonDReg_21),
	.datab(writedata_21),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[21]~17_combout ),
	.cout());
defparam \ociram_wr_data[21]~17 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[21]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[30]~18 (
	.dataa(MonDReg_30),
	.datab(writedata_30),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[30]~18_combout ),
	.cout());
defparam \ociram_wr_data[30]~18 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[30]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[3]~3 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[3]~3_combout ),
	.cout());
defparam \ociram_byteenable[3]~3 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[29]~19 (
	.dataa(MonDReg_29),
	.datab(writedata_29),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[29]~19_combout ),
	.cout());
defparam \ociram_wr_data[29]~19 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[29]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[28]~20 (
	.dataa(MonDReg_28),
	.datab(writedata_28),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[28]~20_combout ),
	.cout());
defparam \ociram_wr_data[28]~20 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[28]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[27]~21 (
	.dataa(MonDReg_27),
	.datab(writedata_27),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[27]~21_combout ),
	.cout());
defparam \ociram_wr_data[27]~21 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[27]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[26]~22 (
	.dataa(MonDReg_26),
	.datab(writedata_26),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[26]~22_combout ),
	.cout());
defparam \ociram_wr_data[26]~22 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[26]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[25]~23 (
	.dataa(MonDReg_25),
	.datab(writedata_25),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[25]~23_combout ),
	.cout());
defparam \ociram_wr_data[25]~23 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[25]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[24]~24 (
	.dataa(MonDReg_24),
	.datab(writedata_24),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[24]~24_combout ),
	.cout());
defparam \ociram_wr_data[24]~24 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[24]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[23]~25 (
	.dataa(MonDReg_23),
	.datab(writedata_23),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[23]~25_combout ),
	.cout());
defparam \ociram_wr_data[23]~25 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[23]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[22]~26 (
	.dataa(MonDReg_22),
	.datab(writedata_22),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[22]~26_combout ),
	.cout());
defparam \ociram_wr_data[22]~26 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[22]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[20]~27 (
	.dataa(MonDReg_20),
	.datab(writedata_20),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[20]~27_combout ),
	.cout());
defparam \ociram_wr_data[20]~27 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[20]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[19]~28 (
	.dataa(MonDReg_19),
	.datab(writedata_19),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[19]~28_combout ),
	.cout());
defparam \ociram_wr_data[19]~28 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[19]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[18]~29 (
	.dataa(MonDReg_18),
	.datab(writedata_18),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[18]~29_combout ),
	.cout());
defparam \ociram_wr_data[18]~29 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[18]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[17]~30 (
	.dataa(MonDReg_17),
	.datab(writedata_17),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[17]~30_combout ),
	.cout());
defparam \ociram_wr_data[17]~30 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[17]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[31]~31 (
	.dataa(MonDReg_31),
	.datab(writedata_31),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[31]~31_combout ),
	.cout());
defparam \ociram_wr_data[31]~31 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[31]~31 .sum_lutc_input = "datac";

dffeas \MonDReg[0] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[0]~0_combout ),
	.asdata(jdo_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[1] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[1]~1_combout ),
	.asdata(jdo_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[3]~2_combout ),
	.asdata(jdo_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[4]~3_combout ),
	.asdata(jdo_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[25]~5_combout ),
	.asdata(jdo_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[26]~4_combout ),
	.asdata(jdo_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[5]~6_combout ),
	.asdata(jdo_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[29]~7_combout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[11]~8_combout ),
	.asdata(jdo_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[12]~9_combout ),
	.asdata(jdo_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[9]~10_combout ),
	.asdata(jdo_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[8]~11_combout ),
	.asdata(jdo_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(take_no_action_ocimem_a),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg[18]~12_combout ),
	.asdata(jdo_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas waitrequest(
	.clk(wire_pll7_clk_0),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[2] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

cycloneive_lcell_comb \ociram_wr_en~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(ociram_wr_en),
	.cout());
defparam \ociram_wr_en~0 .lut_mask = 16'hEEEE;
defparam \ociram_wr_en~0 .sum_lutc_input = "datac";

dffeas \MonDReg[27] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(wire_pll7_clk_0),
	.d(\MonDReg~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~13_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\MonARegAddrInc[0]~0_combout ),
	.cout(\MonARegAddrInc[0]~1 ));
defparam \MonARegAddrInc[0]~0 .lut_mask = 16'h55AA;
defparam \MonARegAddrInc[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonAReg~0 (
	.dataa(jdo_26),
	.datab(\MonARegAddrInc[0]~0_combout ),
	.datac(take_no_action_ocimem_a),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~0_combout ),
	.cout());
defparam \MonAReg~0 .lut_mask = 16'hEFFE;
defparam \MonAReg~0 .sum_lutc_input = "datac";

dffeas \MonAReg[2] (
	.clk(wire_pll7_clk_0),
	.d(\MonAReg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[1]~2 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[0]~1 ),
	.combout(\MonARegAddrInc[1]~2_combout ),
	.cout(\MonARegAddrInc[1]~3 ));
defparam \MonARegAddrInc[1]~2 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~2 (
	.dataa(jdo_27),
	.datab(\MonARegAddrInc[1]~2_combout ),
	.datac(take_no_action_ocimem_a),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~2_combout ),
	.cout());
defparam \MonAReg~2 .lut_mask = 16'hEFFE;
defparam \MonAReg~2 .sum_lutc_input = "datac";

dffeas \MonAReg[3] (
	.clk(wire_pll7_clk_0),
	.d(\MonAReg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[2]~4 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[1]~3 ),
	.combout(\MonARegAddrInc[2]~4_combout ),
	.cout(\MonARegAddrInc[2]~5 ));
defparam \MonARegAddrInc[2]~4 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[2]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~1 (
	.dataa(jdo_28),
	.datab(\MonARegAddrInc[2]~4_combout ),
	.datac(take_no_action_ocimem_a),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~1_combout ),
	.cout());
defparam \MonAReg~1 .lut_mask = 16'hEFFE;
defparam \MonAReg~1 .sum_lutc_input = "datac";

dffeas \MonAReg[4] (
	.clk(wire_pll7_clk_0),
	.d(\MonAReg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hAFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_access~0 (
	.dataa(jdo_17),
	.datab(\MonARegAddrInc[8]~16_combout ),
	.datac(take_no_action_ocimem_a),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.cout());
defparam \jtag_ram_access~0 .lut_mask = 16'hEFFE;
defparam \jtag_ram_access~0 .sum_lutc_input = "datac";

dffeas \MonAReg[10] (
	.clk(wire_pll7_clk_0),
	.d(\jtag_ram_access~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[3]~6 (
	.dataa(\MonAReg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[2]~5 ),
	.combout(\MonARegAddrInc[3]~6_combout ),
	.cout(\MonARegAddrInc[3]~7 ));
defparam \MonARegAddrInc[3]~6 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~3 (
	.dataa(jdo_29),
	.datab(\MonARegAddrInc[3]~6_combout ),
	.datac(take_no_action_ocimem_a),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~3_combout ),
	.cout());
defparam \MonAReg~3 .lut_mask = 16'hEFFE;
defparam \MonAReg~3 .sum_lutc_input = "datac";

dffeas \MonAReg[5] (
	.clk(wire_pll7_clk_0),
	.d(\MonAReg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[4]~8 (
	.dataa(\MonAReg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[3]~7 ),
	.combout(\MonARegAddrInc[4]~8_combout ),
	.cout(\MonARegAddrInc[4]~9 ));
defparam \MonARegAddrInc[4]~8 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[4]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~4 (
	.dataa(jdo_30),
	.datab(\MonARegAddrInc[4]~8_combout ),
	.datac(take_no_action_ocimem_a),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~4_combout ),
	.cout());
defparam \MonAReg~4 .lut_mask = 16'hEFFE;
defparam \MonAReg~4 .sum_lutc_input = "datac";

dffeas \MonAReg[6] (
	.clk(wire_pll7_clk_0),
	.d(\MonAReg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[5]~10 (
	.dataa(\MonAReg[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[4]~9 ),
	.combout(\MonARegAddrInc[5]~10_combout ),
	.cout(\MonARegAddrInc[5]~11 ));
defparam \MonARegAddrInc[5]~10 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[5]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~5 (
	.dataa(jdo_31),
	.datab(\MonARegAddrInc[5]~10_combout ),
	.datac(take_no_action_ocimem_a),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~5_combout ),
	.cout());
defparam \MonAReg~5 .lut_mask = 16'hEFFE;
defparam \MonAReg~5 .sum_lutc_input = "datac";

dffeas \MonAReg[7] (
	.clk(wire_pll7_clk_0),
	.d(\MonAReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[6]~12 (
	.dataa(\MonAReg[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[5]~11 ),
	.combout(\MonARegAddrInc[6]~12_combout ),
	.cout(\MonARegAddrInc[6]~13 ));
defparam \MonARegAddrInc[6]~12 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[6]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~6 (
	.dataa(jdo_32),
	.datab(\MonARegAddrInc[6]~12_combout ),
	.datac(take_no_action_ocimem_a),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~6_combout ),
	.cout());
defparam \MonAReg~6 .lut_mask = 16'hEFFE;
defparam \MonAReg~6 .sum_lutc_input = "datac";

dffeas \MonAReg[8] (
	.clk(wire_pll7_clk_0),
	.d(\MonAReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[7]~14 (
	.dataa(\MonAReg[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[6]~13 ),
	.combout(\MonARegAddrInc[7]~14_combout ),
	.cout(\MonARegAddrInc[7]~15 ));
defparam \MonARegAddrInc[7]~14 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[7]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~7 (
	.dataa(jdo_33),
	.datab(\MonARegAddrInc[7]~14_combout ),
	.datac(take_no_action_ocimem_a),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~7_combout ),
	.cout());
defparam \MonAReg~7 .lut_mask = 16'hEFFE;
defparam \MonAReg~7 .sum_lutc_input = "datac";

dffeas \MonAReg[9] (
	.clk(wire_pll7_clk_0),
	.d(\MonAReg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[8]~16 (
	.dataa(\MonAReg[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\MonARegAddrInc[7]~15 ),
	.combout(\MonARegAddrInc[8]~16_combout ),
	.cout());
defparam \MonARegAddrInc[8]~16 .lut_mask = 16'h5A5A;
defparam \MonARegAddrInc[8]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \jtag_ram_rd~0 (
	.dataa(take_no_action_ocimem_a),
	.datab(jdo_34),
	.datac(\MonARegAddrInc[8]~16_combout ),
	.datad(jdo_17),
	.cin(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.cout());
defparam \jtag_ram_rd~0 .lut_mask = 16'h47FF;
defparam \jtag_ram_rd~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_rd~1 (
	.dataa(\jtag_ram_rd~0_combout ),
	.datab(take_action_ocimem_b),
	.datac(\jtag_ram_rd~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\jtag_ram_rd~1_combout ),
	.cout());
defparam \jtag_ram_rd~1 .lut_mask = 16'hFEFE;
defparam \jtag_ram_rd~1 .sum_lutc_input = "datac";

dffeas jtag_ram_rd(
	.clk(wire_pll7_clk_0),
	.d(\jtag_ram_rd~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(wire_pll7_clk_0),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cycloneive_lcell_comb \MonDReg[0]~0 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_0),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[0]~0_combout ),
	.cout());
defparam \MonDReg[0]~0 .lut_mask = 16'hAACC;
defparam \MonDReg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_rd~0 (
	.dataa(take_action_ocimem_a),
	.datab(\jtag_rd~q ),
	.datac(gnd),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\jtag_rd~0_combout ),
	.cout());
defparam \jtag_rd~0 .lut_mask = 16'hEEFF;
defparam \jtag_rd~0 .sum_lutc_input = "datac";

dffeas jtag_rd(
	.clk(wire_pll7_clk_0),
	.d(\jtag_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(wire_pll7_clk_0),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cycloneive_lcell_comb \MonDReg[0]~13 (
	.dataa(take_no_action_ocimem_a),
	.datab(gnd),
	.datac(take_action_ocimem_b),
	.datad(\jtag_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[0]~13_combout ),
	.cout());
defparam \MonDReg[0]~13 .lut_mask = 16'hFFFA;
defparam \MonDReg[0]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[1]~1 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_1),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[1]~1_combout ),
	.cout());
defparam \MonDReg[1]~1 .lut_mask = 16'hAACC;
defparam \MonDReg[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[3]~2 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_3),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[3]~2_combout ),
	.cout());
defparam \MonDReg[3]~2 .lut_mask = 16'hAACC;
defparam \MonDReg[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[4]~3 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_4),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[4]~3_combout ),
	.cout());
defparam \MonDReg[4]~3 .lut_mask = 16'hAACC;
defparam \MonDReg[4]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(gnd),
	.datab(\MonAReg[4]~q ),
	.datac(\MonAReg[3]~q ),
	.datad(\MonAReg[2]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h3FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[25]~5 (
	.dataa(\Equal0~1_combout ),
	.datab(q_a_25),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[25]~5_combout ),
	.cout());
defparam \MonDReg[25]~5 .lut_mask = 16'hAACC;
defparam \MonDReg[25]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\MonAReg[4]~q ),
	.datab(\MonAReg[2]~q ),
	.datac(gnd),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[26]~4 (
	.dataa(\Equal0~2_combout ),
	.datab(q_a_26),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[26]~4_combout ),
	.cout());
defparam \MonDReg[26]~4 .lut_mask = 16'hAACC;
defparam \MonDReg[26]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[5]~6 (
	.dataa(\Equal0~1_combout ),
	.datab(q_a_5),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[5]~6_combout ),
	.cout());
defparam \MonDReg[5]~6 .lut_mask = 16'hAACC;
defparam \MonDReg[5]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(\MonAReg[3]~q ),
	.datad(\MonAReg[2]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hAFFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[29]~7 (
	.dataa(\Equal0~3_combout ),
	.datab(q_a_29),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[29]~7_combout ),
	.cout());
defparam \MonDReg[29]~7 .lut_mask = 16'hAACC;
defparam \MonDReg[29]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[11]~8 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_11),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[11]~8_combout ),
	.cout());
defparam \MonDReg[11]~8 .lut_mask = 16'hAACC;
defparam \MonDReg[11]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'hAAFF;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[12]~9 (
	.dataa(\Equal0~4_combout ),
	.datab(q_a_12),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[12]~9_combout ),
	.cout());
defparam \MonDReg[12]~9 .lut_mask = 16'hAACC;
defparam \MonDReg[12]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[9]~10 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_9),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[9]~10_combout ),
	.cout());
defparam \MonDReg[9]~10 .lut_mask = 16'hAACC;
defparam \MonDReg[9]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~28 (
	.dataa(q_a_8),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\MonDReg~28_combout ),
	.cout());
defparam \MonDReg~28 .lut_mask = 16'hB8FF;
defparam \MonDReg~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[8]~11 (
	.dataa(MonDReg_8),
	.datab(\MonDReg~28_combout ),
	.datac(gnd),
	.datad(\jtag_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[8]~11_combout ),
	.cout());
defparam \MonDReg[8]~11 .lut_mask = 16'hAACC;
defparam \MonDReg[8]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~5 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[2]~q ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'hAFFF;
defparam \Equal0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[18]~12 (
	.dataa(\Equal0~5_combout ),
	.datab(q_a_18),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[18]~12_combout ),
	.cout());
defparam \MonDReg[18]~12 .lut_mask = 16'hAACC;
defparam \MonDReg[18]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_access~1 (
	.dataa(\jtag_ram_access~0_combout ),
	.datab(\MonARegAddrInc[8]~16_combout ),
	.datac(take_action_ocimem_b),
	.datad(take_no_action_ocimem_a),
	.cin(gnd),
	.combout(\jtag_ram_access~1_combout ),
	.cout());
defparam \jtag_ram_access~1 .lut_mask = 16'hF377;
defparam \jtag_ram_access~1 .sum_lutc_input = "datac";

dffeas jtag_ram_access(
	.clk(wire_pll7_clk_0),
	.d(\jtag_ram_access~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cycloneive_lcell_comb \waitrequest~0 (
	.dataa(write),
	.datab(\jtag_ram_access~q ),
	.datac(address_8),
	.datad(waitrequest1),
	.cin(gnd),
	.combout(\waitrequest~0_combout ),
	.cout());
defparam \waitrequest~0 .lut_mask = 16'hEFFF;
defparam \waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(read),
	.datab(address_8),
	.datac(\jtag_ram_access~q ),
	.datad(write),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 16'hEFFF;
defparam \avalon_ociram_readdata_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avalon_ociram_readdata_ready~1 (
	.dataa(waitrequest1),
	.datab(\avalon_ociram_readdata_ready~0_combout ),
	.datac(write),
	.datad(\avalon_ociram_readdata_ready~q ),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~1_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~1 .lut_mask = 16'hFFFE;
defparam \avalon_ociram_readdata_ready~1 .sum_lutc_input = "datac";

dffeas avalon_ociram_readdata_ready(
	.clk(wire_pll7_clk_0),
	.d(\avalon_ociram_readdata_ready~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cycloneive_lcell_comb \waitrequest~1 (
	.dataa(\waitrequest~0_combout ),
	.datab(read),
	.datac(\avalon_ociram_readdata_ready~q ),
	.datad(write),
	.cin(gnd),
	.combout(\waitrequest~1_combout ),
	.cout());
defparam \waitrequest~1 .lut_mask = 16'hBFFF;
defparam \waitrequest~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~14 (
	.dataa(jdo_5),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_2),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~14_combout ),
	.cout());
defparam \MonDReg~14 .lut_mask = 16'hFAFC;
defparam \MonDReg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~15 (
	.dataa(jdo_30),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_27),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~15_combout ),
	.cout());
defparam \MonDReg~15 .lut_mask = 16'hFAFC;
defparam \MonDReg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~16 (
	.dataa(jdo_27),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_24),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~16_combout ),
	.cout());
defparam \MonDReg~16 .lut_mask = 16'hFAFC;
defparam \MonDReg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~17 (
	.dataa(jdo_19),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_16),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~17_combout ),
	.cout());
defparam \MonDReg~17 .lut_mask = 16'hFAFC;
defparam \MonDReg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~18 (
	.dataa(jdo_23),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_20),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~18_combout ),
	.cout());
defparam \MonDReg~18 .lut_mask = 16'hFAFC;
defparam \MonDReg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~19 (
	.dataa(jdo_22),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_19),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~19_combout ),
	.cout());
defparam \MonDReg~19 .lut_mask = 16'hFAFC;
defparam \MonDReg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~20 (
	.dataa(jdo_31),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_28),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~20_combout ),
	.cout());
defparam \MonDReg~20 .lut_mask = 16'hFAFC;
defparam \MonDReg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~21 (
	.dataa(jdo_33),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_30),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~21_combout ),
	.cout());
defparam \MonDReg~21 .lut_mask = 16'hFAFC;
defparam \MonDReg~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~22 (
	.dataa(jdo_34),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_31),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~22_combout ),
	.cout());
defparam \MonDReg~22 .lut_mask = 16'hFAFC;
defparam \MonDReg~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~23 (
	.dataa(jdo_20),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_17),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~23_combout ),
	.cout());
defparam \MonDReg~23 .lut_mask = 16'hFAFC;
defparam \MonDReg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~24 (
	.dataa(jdo_16),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_13),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~24_combout ),
	.cout());
defparam \MonDReg~24 .lut_mask = 16'hFAFC;
defparam \MonDReg~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~25 (
	.dataa(jdo_17),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_14),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~25_combout ),
	.cout());
defparam \MonDReg~25 .lut_mask = 16'hFAFC;
defparam \MonDReg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~26 (
	.dataa(jdo_18),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_15),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~26_combout ),
	.cout());
defparam \MonDReg~26 .lut_mask = 16'hFAFC;
defparam \MonDReg~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~27 (
	.dataa(jdo_13),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_10),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~27_combout ),
	.cout());
defparam \MonDReg~27 .lut_mask = 16'hFAFC;
defparam \MonDReg~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~29 (
	.dataa(jdo_10),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_7),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~29_combout ),
	.cout());
defparam \MonDReg~29 .lut_mask = 16'hFAFC;
defparam \MonDReg~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~30 (
	.dataa(jdo_9),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_6),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~30_combout ),
	.cout());
defparam \MonDReg~30 .lut_mask = 16'hFAFC;
defparam \MonDReg~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~31 (
	.dataa(jdo_24),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_21),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~31_combout ),
	.cout());
defparam \MonDReg~31 .lut_mask = 16'hFAFC;
defparam \MonDReg~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~32 (
	.dataa(jdo_26),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_23),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~32_combout ),
	.cout());
defparam \MonDReg~32 .lut_mask = 16'hFAFC;
defparam \MonDReg~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~33 (
	.dataa(jdo_25),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_22),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~33_combout ),
	.cout());
defparam \MonDReg~33 .lut_mask = 16'hFAFC;
defparam \MonDReg~33 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_cpu_cpu_ociram_sp_ram_module (
	wire_pll7_clk_0,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_21,
	q_a_30,
	q_a_29,
	q_a_28,
	q_a_27,
	q_a_26,
	q_a_25,
	q_a_24,
	q_a_23,
	q_a_22,
	q_a_20,
	q_a_19,
	q_a_18,
	q_a_17,
	q_a_31,
	ociram_wr_en,
	ociram_reset_req,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_3,
	ociram_wr_data_4,
	ociram_wr_data_11,
	ociram_byteenable_1,
	ociram_wr_data_13,
	ociram_wr_data_16,
	ociram_byteenable_2,
	ociram_wr_data_12,
	ociram_wr_data_5,
	ociram_wr_data_14,
	ociram_wr_data_15,
	ociram_wr_data_10,
	ociram_wr_data_9,
	ociram_wr_data_8,
	ociram_wr_data_7,
	ociram_wr_data_6,
	ociram_wr_data_21,
	ociram_wr_data_30,
	ociram_byteenable_3,
	ociram_wr_data_29,
	ociram_wr_data_28,
	ociram_wr_data_27,
	ociram_wr_data_26,
	ociram_wr_data_25,
	ociram_wr_data_24,
	ociram_wr_data_23,
	ociram_wr_data_22,
	ociram_wr_data_20,
	ociram_wr_data_19,
	ociram_wr_data_18,
	ociram_wr_data_17,
	ociram_wr_data_31)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_10;
output 	q_a_9;
output 	q_a_8;
output 	q_a_7;
output 	q_a_6;
output 	q_a_21;
output 	q_a_30;
output 	q_a_29;
output 	q_a_28;
output 	q_a_27;
output 	q_a_26;
output 	q_a_25;
output 	q_a_24;
output 	q_a_23;
output 	q_a_22;
output 	q_a_20;
output 	q_a_19;
output 	q_a_18;
output 	q_a_17;
output 	q_a_31;
input 	ociram_wr_en;
input 	ociram_reset_req;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_3;
input 	ociram_wr_data_4;
input 	ociram_wr_data_11;
input 	ociram_byteenable_1;
input 	ociram_wr_data_13;
input 	ociram_wr_data_16;
input 	ociram_byteenable_2;
input 	ociram_wr_data_12;
input 	ociram_wr_data_5;
input 	ociram_wr_data_14;
input 	ociram_wr_data_15;
input 	ociram_wr_data_10;
input 	ociram_wr_data_9;
input 	ociram_wr_data_8;
input 	ociram_wr_data_7;
input 	ociram_wr_data_6;
input 	ociram_wr_data_21;
input 	ociram_wr_data_30;
input 	ociram_byteenable_3;
input 	ociram_wr_data_29;
input 	ociram_wr_data_28;
input 	ociram_wr_data_27;
input 	ociram_wr_data_26;
input 	ociram_wr_data_25;
input 	ociram_wr_data_24;
input 	ociram_wr_data_23;
input 	ociram_wr_data_22;
input 	ociram_wr_data_20;
input 	ociram_wr_data_19;
input 	ociram_wr_data_18;
input 	ociram_wr_data_17;
input 	ociram_wr_data_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altsyncram_1 the_altsyncram(
	.clock0(wire_pll7_clk_0),
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(ociram_reset_req),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}));

endmodule

module niosII_altsyncram_1 (
	clock0,
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altsyncram_ac71 auto_generated(
	.clock0(clock0),
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}));

endmodule

module niosII_altsyncram_ac71 (
	clock0,
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_nios2_oci:the_niosII_cpu_cpu_nios2_oci|niosII_cpu_cpu_nios2_ocimem:the_niosII_cpu_cpu_nios2_ocimem|niosII_cpu_cpu_ociram_sp_ram_module:niosII_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module niosII_niosII_cpu_cpu_register_bank_a_module (
	wire_pll7_clk_0,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_31,
	q_b_30,
	q_b_29,
	q_b_28,
	q_b_27,
	D_iw_30,
	D_iw_29,
	D_iw_28,
	D_iw_27,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	D_iw_31,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_24,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	W_rf_wr_data_16,
	W_rf_wr_data_15,
	W_rf_wr_data_14,
	W_rf_wr_data_13,
	W_rf_wr_data_12,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_9,
	W_rf_wr_data_8,
	W_rf_wr_data_27,
	W_rf_wr_data_28,
	W_rf_wr_data_29,
	W_rf_wr_data_30,
	W_rf_wr_data_31)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
output 	q_b_28;
output 	q_b_27;
input 	D_iw_30;
input 	D_iw_29;
input 	D_iw_28;
input 	D_iw_27;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	D_iw_31;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_29;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altsyncram_2 the_altsyncram(
	.clock0(wire_pll7_clk_0),
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({D_iw_31,D_iw_30,D_iw_29,D_iw_28,D_iw_27}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}));

endmodule

module niosII_altsyncram_2 (
	clock0,
	q_b,
	address_b,
	wren_a,
	data_a,
	address_a)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altsyncram_6mc1 auto_generated(
	.clock0(clock0),
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}));

endmodule

module niosII_altsyncram_6mc1 (
	clock0,
	q_b,
	address_b,
	wren_a,
	data_a,
	address_a)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_a_module:niosII_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

endmodule

module niosII_niosII_cpu_cpu_register_bank_b_module (
	wire_pll7_clk_0,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	D_iw_26,
	D_iw_25,
	D_iw_24,
	D_iw_23,
	D_iw_22,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_24,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	W_rf_wr_data_16,
	W_rf_wr_data_15,
	W_rf_wr_data_14,
	W_rf_wr_data_13,
	W_rf_wr_data_12,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_9,
	W_rf_wr_data_8,
	W_rf_wr_data_27,
	W_rf_wr_data_28,
	W_rf_wr_data_29,
	W_rf_wr_data_30,
	W_rf_wr_data_31)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
input 	D_iw_26;
input 	D_iw_25;
input 	D_iw_24;
input 	D_iw_23;
input 	D_iw_22;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_29;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altsyncram_3 the_altsyncram(
	.clock0(wire_pll7_clk_0),
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({D_iw_26,D_iw_25,D_iw_24,D_iw_23,D_iw_22}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}));

endmodule

module niosII_altsyncram_3 (
	clock0,
	q_b,
	address_b,
	wren_a,
	data_a,
	address_a)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altsyncram_6mc1_1 auto_generated(
	.clock0(clock0),
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}));

endmodule

module niosII_altsyncram_6mc1_1 (
	clock0,
	q_b,
	address_b,
	wren_a,
	data_a,
	address_a)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "niosII_cpu:cpu|niosII_cpu_cpu:cpu|niosII_cpu_cpu_register_bank_b_module:niosII_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module niosII_niosII_epcs (
	wire_pll7_clk_0,
	SCLK_reg,
	sce,
	shift_reg_7,
	r_sync_rst,
	saved_grant_0,
	saved_grant_1,
	out_data_buffer_38,
	src_data_38,
	src_data_39,
	src_data_40,
	src_payload,
	src_payload1,
	mem_used_1,
	wait_latency_counter_1,
	src_valid,
	src_valid1,
	src_data_46,
	out_data_buffer_65,
	p1_wr_strobe,
	src_payload2,
	src_payload3,
	src_data_66,
	av_begintransfer,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_14,
	readdata_15,
	readdata_10,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_6,
	readdata_21,
	readdata_30,
	readdata_29,
	readdata_28,
	readdata_27,
	readdata_26,
	readdata_25,
	readdata_24,
	readdata_23,
	readdata_22,
	readdata_20,
	readdata_19,
	readdata_18,
	readdata_17,
	src_payload9,
	irq_reg,
	r_early_rst,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_payload10,
	readdata_31,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	epcs_data0)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	SCLK_reg;
output 	sce;
output 	shift_reg_7;
input 	r_sync_rst;
input 	saved_grant_0;
input 	saved_grant_1;
input 	out_data_buffer_38;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_payload;
input 	src_payload1;
input 	mem_used_1;
input 	wait_latency_counter_1;
input 	src_valid;
input 	src_valid1;
input 	src_data_46;
input 	out_data_buffer_65;
output 	p1_wr_strobe;
input 	src_payload2;
input 	src_payload3;
input 	src_data_66;
input 	av_begintransfer;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_5;
output 	readdata_14;
output 	readdata_15;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_6;
output 	readdata_21;
output 	readdata_30;
output 	readdata_29;
output 	readdata_28;
output 	readdata_27;
output 	readdata_26;
output 	readdata_25;
output 	readdata_24;
output 	readdata_23;
output 	readdata_22;
output 	readdata_20;
output 	readdata_19;
output 	readdata_18;
output 	readdata_17;
input 	src_payload9;
output 	irq_reg;
input 	r_early_rst;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_payload10;
output 	readdata_31;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	epcs_data0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_boot_copier_rom|auto_generated|q_a[0] ;
wire \the_boot_copier_rom|auto_generated|q_a[1] ;
wire \the_boot_copier_rom|auto_generated|q_a[2] ;
wire \the_boot_copier_rom|auto_generated|q_a[3] ;
wire \the_boot_copier_rom|auto_generated|q_a[4] ;
wire \the_boot_copier_rom|auto_generated|q_a[11] ;
wire \the_boot_copier_rom|auto_generated|q_a[13] ;
wire \the_boot_copier_rom|auto_generated|q_a[16] ;
wire \the_boot_copier_rom|auto_generated|q_a[12] ;
wire \the_niosII_epcs_sub|data_to_cpu[5]~q ;
wire \the_boot_copier_rom|auto_generated|q_a[5] ;
wire \the_boot_copier_rom|auto_generated|q_a[14] ;
wire \the_boot_copier_rom|auto_generated|q_a[15] ;
wire \the_boot_copier_rom|auto_generated|q_a[10] ;
wire \the_boot_copier_rom|auto_generated|q_a[9] ;
wire \the_boot_copier_rom|auto_generated|q_a[8] ;
wire \the_boot_copier_rom|auto_generated|q_a[7] ;
wire \the_boot_copier_rom|auto_generated|q_a[6] ;
wire \the_boot_copier_rom|auto_generated|q_a[21] ;
wire \the_boot_copier_rom|auto_generated|q_a[30] ;
wire \the_boot_copier_rom|auto_generated|q_a[29] ;
wire \the_boot_copier_rom|auto_generated|q_a[28] ;
wire \the_boot_copier_rom|auto_generated|q_a[27] ;
wire \the_boot_copier_rom|auto_generated|q_a[26] ;
wire \the_boot_copier_rom|auto_generated|q_a[25] ;
wire \the_boot_copier_rom|auto_generated|q_a[24] ;
wire \the_boot_copier_rom|auto_generated|q_a[23] ;
wire \the_boot_copier_rom|auto_generated|q_a[22] ;
wire \the_boot_copier_rom|auto_generated|q_a[20] ;
wire \the_boot_copier_rom|auto_generated|q_a[19] ;
wire \the_boot_copier_rom|auto_generated|q_a[18] ;
wire \the_boot_copier_rom|auto_generated|q_a[17] ;
wire \the_boot_copier_rom|auto_generated|q_a[31] ;
wire \the_niosII_epcs_sub|data_to_cpu[0]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[1]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[2]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[3]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[4]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[11]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[13]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[12]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[14]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[15]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[10]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[9]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[8]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[7]~q ;
wire \the_niosII_epcs_sub|data_to_cpu[6]~q ;


niosII_altsyncram_4 the_boot_copier_rom(
	.clock0(wire_pll7_clk_0),
	.q_a({\the_boot_copier_rom|auto_generated|q_a[31] ,\the_boot_copier_rom|auto_generated|q_a[30] ,\the_boot_copier_rom|auto_generated|q_a[29] ,\the_boot_copier_rom|auto_generated|q_a[28] ,\the_boot_copier_rom|auto_generated|q_a[27] ,
\the_boot_copier_rom|auto_generated|q_a[26] ,\the_boot_copier_rom|auto_generated|q_a[25] ,\the_boot_copier_rom|auto_generated|q_a[24] ,\the_boot_copier_rom|auto_generated|q_a[23] ,\the_boot_copier_rom|auto_generated|q_a[22] ,
\the_boot_copier_rom|auto_generated|q_a[21] ,\the_boot_copier_rom|auto_generated|q_a[20] ,\the_boot_copier_rom|auto_generated|q_a[19] ,\the_boot_copier_rom|auto_generated|q_a[18] ,\the_boot_copier_rom|auto_generated|q_a[17] ,
\the_boot_copier_rom|auto_generated|q_a[16] ,\the_boot_copier_rom|auto_generated|q_a[15] ,\the_boot_copier_rom|auto_generated|q_a[14] ,\the_boot_copier_rom|auto_generated|q_a[13] ,\the_boot_copier_rom|auto_generated|q_a[12] ,
\the_boot_copier_rom|auto_generated|q_a[11] ,\the_boot_copier_rom|auto_generated|q_a[10] ,\the_boot_copier_rom|auto_generated|q_a[9] ,\the_boot_copier_rom|auto_generated|q_a[8] ,\the_boot_copier_rom|auto_generated|q_a[7] ,
\the_boot_copier_rom|auto_generated|q_a[6] ,\the_boot_copier_rom|auto_generated|q_a[5] ,\the_boot_copier_rom|auto_generated|q_a[4] ,\the_boot_copier_rom|auto_generated|q_a[3] ,\the_boot_copier_rom|auto_generated|q_a[2] ,
\the_boot_copier_rom|auto_generated|q_a[1] ,\the_boot_copier_rom|auto_generated|q_a[0] }),
	.address_a({src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.clocken0(r_early_rst));

niosII_niosII_epcs_sub the_niosII_epcs_sub(
	.clk(wire_pll7_clk_0),
	.data_to_cpu_5(\the_niosII_epcs_sub|data_to_cpu[5]~q ),
	.SCLK_reg1(SCLK_reg),
	.SS_n(sce),
	.shift_reg_7(shift_reg_7),
	.reset_n(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.saved_grant_1(saved_grant_1),
	.out_data_buffer_38(out_data_buffer_38),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.data_from_cpu({src_payload15,src_payload14,src_payload12,src_payload13,src_payload11,src_payload,src_payload16,src_payload17,src_payload2,src_payload4,src_payload5,src_payload6,src_payload7,src_payload8,src_payload9,src_payload1}),
	.mem_used_1(mem_used_1),
	.wait_latency_counter_1(wait_latency_counter_1),
	.src_valid(src_valid),
	.src_valid1(src_valid1),
	.src_data_46(src_data_46),
	.out_data_buffer_65(out_data_buffer_65),
	.p1_wr_strobe(p1_wr_strobe),
	.src_payload(src_payload3),
	.src_data_66(src_data_66),
	.data_to_cpu_0(\the_niosII_epcs_sub|data_to_cpu[0]~q ),
	.data_to_cpu_1(\the_niosII_epcs_sub|data_to_cpu[1]~q ),
	.data_to_cpu_2(\the_niosII_epcs_sub|data_to_cpu[2]~q ),
	.data_to_cpu_3(\the_niosII_epcs_sub|data_to_cpu[3]~q ),
	.data_to_cpu_4(\the_niosII_epcs_sub|data_to_cpu[4]~q ),
	.data_to_cpu_11(\the_niosII_epcs_sub|data_to_cpu[11]~q ),
	.data_to_cpu_13(\the_niosII_epcs_sub|data_to_cpu[13]~q ),
	.data_to_cpu_12(\the_niosII_epcs_sub|data_to_cpu[12]~q ),
	.data_to_cpu_14(\the_niosII_epcs_sub|data_to_cpu[14]~q ),
	.data_to_cpu_15(\the_niosII_epcs_sub|data_to_cpu[15]~q ),
	.data_to_cpu_10(\the_niosII_epcs_sub|data_to_cpu[10]~q ),
	.data_to_cpu_9(\the_niosII_epcs_sub|data_to_cpu[9]~q ),
	.data_to_cpu_8(\the_niosII_epcs_sub|data_to_cpu[8]~q ),
	.data_to_cpu_7(\the_niosII_epcs_sub|data_to_cpu[7]~q ),
	.data_to_cpu_6(\the_niosII_epcs_sub|data_to_cpu[6]~q ),
	.irq_reg1(irq_reg),
	.src_payload1(src_payload10),
	.epcs_data0(epcs_data0));

cycloneive_lcell_comb \readdata[0]~0 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[0]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[0] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0]~0 .lut_mask = 16'hEFFE;
defparam \readdata[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1]~1 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[1]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[1] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1]~1 .lut_mask = 16'hEFFE;
defparam \readdata[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[2]~2 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[2]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[2] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2]~2 .lut_mask = 16'hEFFE;
defparam \readdata[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3]~3 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[3]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[3] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3]~3 .lut_mask = 16'hEFFE;
defparam \readdata[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[4]~4 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[4]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[4] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4]~4 .lut_mask = 16'hEFFE;
defparam \readdata[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[11]~5 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[11]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[11] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_11),
	.cout());
defparam \readdata[11]~5 .lut_mask = 16'hEFFE;
defparam \readdata[11]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[13]~6 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[13]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[13] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_13),
	.cout());
defparam \readdata[13]~6 .lut_mask = 16'hEFFE;
defparam \readdata[13]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[16]~7 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[16] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_16),
	.cout());
defparam \readdata[16]~7 .lut_mask = 16'hAFFF;
defparam \readdata[16]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[12]~8 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[12]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[12] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_12),
	.cout());
defparam \readdata[12]~8 .lut_mask = 16'hEFFE;
defparam \readdata[12]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[5]~9 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[5]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[5] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5]~9 .lut_mask = 16'hEFFE;
defparam \readdata[5]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[14]~10 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[14]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[14] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_14),
	.cout());
defparam \readdata[14]~10 .lut_mask = 16'hEFFE;
defparam \readdata[14]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[15]~11 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[15]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[15] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_15),
	.cout());
defparam \readdata[15]~11 .lut_mask = 16'hEFFE;
defparam \readdata[15]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[10]~12 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[10]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[10] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_10),
	.cout());
defparam \readdata[10]~12 .lut_mask = 16'hEFFE;
defparam \readdata[10]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[9]~13 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[9]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[9] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_9),
	.cout());
defparam \readdata[9]~13 .lut_mask = 16'hEFFE;
defparam \readdata[9]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[8]~14 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[8]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[8] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_8),
	.cout());
defparam \readdata[8]~14 .lut_mask = 16'hEFFE;
defparam \readdata[8]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[7]~15 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[7]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[7] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7]~15 .lut_mask = 16'hEFFE;
defparam \readdata[7]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[6]~16 (
	.dataa(\the_niosII_epcs_sub|data_to_cpu[6]~q ),
	.datab(\the_boot_copier_rom|auto_generated|q_a[6] ),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6]~16 .lut_mask = 16'hEFFE;
defparam \readdata[6]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[21]~17 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[21] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_21),
	.cout());
defparam \readdata[21]~17 .lut_mask = 16'hAFFF;
defparam \readdata[21]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[30]~18 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[30] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_30),
	.cout());
defparam \readdata[30]~18 .lut_mask = 16'hAFFF;
defparam \readdata[30]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[29]~19 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[29] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_29),
	.cout());
defparam \readdata[29]~19 .lut_mask = 16'hAFFF;
defparam \readdata[29]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[28]~20 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[28] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_28),
	.cout());
defparam \readdata[28]~20 .lut_mask = 16'hAFFF;
defparam \readdata[28]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[27]~21 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[27] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_27),
	.cout());
defparam \readdata[27]~21 .lut_mask = 16'hAFFF;
defparam \readdata[27]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[26]~22 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[26] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_26),
	.cout());
defparam \readdata[26]~22 .lut_mask = 16'hAFFF;
defparam \readdata[26]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[25]~23 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[25] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_25),
	.cout());
defparam \readdata[25]~23 .lut_mask = 16'hAFFF;
defparam \readdata[25]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[24]~24 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[24] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_24),
	.cout());
defparam \readdata[24]~24 .lut_mask = 16'hAFFF;
defparam \readdata[24]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[23]~25 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[23] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_23),
	.cout());
defparam \readdata[23]~25 .lut_mask = 16'hAFFF;
defparam \readdata[23]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[22]~26 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[22] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_22),
	.cout());
defparam \readdata[22]~26 .lut_mask = 16'hAFFF;
defparam \readdata[22]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[20]~27 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[20] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_20),
	.cout());
defparam \readdata[20]~27 .lut_mask = 16'hAFFF;
defparam \readdata[20]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[19]~28 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[19] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_19),
	.cout());
defparam \readdata[19]~28 .lut_mask = 16'hAFFF;
defparam \readdata[19]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[18]~29 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[18] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_18),
	.cout());
defparam \readdata[18]~29 .lut_mask = 16'hAFFF;
defparam \readdata[18]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[17]~30 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[17] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_17),
	.cout());
defparam \readdata[17]~30 .lut_mask = 16'hAFFF;
defparam \readdata[17]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[31]~31 (
	.dataa(\the_boot_copier_rom|auto_generated|q_a[31] ),
	.datab(gnd),
	.datac(src_data_46),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(readdata_31),
	.cout());
defparam \readdata[31]~31 .lut_mask = 16'hAFFF;
defparam \readdata[31]~31 .sum_lutc_input = "datac";

endmodule

module niosII_altsyncram_4 (
	clock0,
	q_a,
	address_a,
	clocken0)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_a;
input 	[7:0] address_a;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altsyncram_0941 auto_generated(
	.clock0(clock0),
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clocken0(clocken0));

endmodule

module niosII_altsyncram_0941 (
	clock0,
	q_a,
	address_a,
	clocken0)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_a;
input 	[7:0] address_a;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 256'h00000000000000000000000004C800081228820000211449001064E640000000;

cycloneive_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 256'h000000000001FADDF977E2E62EABBEB6C58629EEDF8AC31577A7B63557FFFEF5;

cycloneive_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 256'h000000000000A763578D5FDDD3FCC94DBF7DFB55A975BEFFCD7C7FFFEEADA59A;

cycloneive_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 256'h00000000000158DEA97AA2A22913B6B2408224AA568A410232838A0891525A75;

cycloneive_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 256'h00000000000158DCA972A2A268CBB6BA52AAA2AA56AB55493A93A66651525A77;

cycloneive_ram_block ram_block1a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "rom";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = 256'h00000000000103E0058D135C4A23C0B405442949130A22162305921134E54D1C;

cycloneive_ram_block ram_block1a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "rom";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = 256'h000000000001F170E9C3A3F26B21D41340C201E10DC2610410829A1927FB3779;

cycloneive_ram_block ram_block1a16(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "rom";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = 256'h000000000000A3E1518543440222C0A00810400A12180824220912113489491D;

cycloneive_ram_block ram_block1a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "rom";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = 256'h000000000000297D41F543104230F200810408010900200411041211A4892599;

cycloneive_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 256'h0000000000015A9CA872A0222EEB36BA52AA8EAED6AB555D3AB3F4F75153DA67;

cycloneive_ram_block ram_block1a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "rom";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = 256'h000000000001FB69E9A7A3626A21C412408200A04482C3044982921125DB375D;

cycloneive_ram_block ram_block1a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "rom";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = 256'h00000000000059FDB9F6E3666222D4A2408200A8568841043A83121135DB5BD8;

cycloneive_ram_block ram_block1a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "rom";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = 256'h000000000000032600951594422068042044240008400014402410112689A190;

cycloneive_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = 256'h00000000000003241095075040886A0C922C86458861B4494414040464812500;

cycloneive_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = 256'h0000000000002520428103145264C14C376DA341816514CCC13410532EA92110;

cycloneive_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 256'h0000000000000D24029001104000400020410001004000800040000020000100;

cycloneive_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 256'h0000000000000D2C06A00510C000400020401411204020000040010020000102;

cycloneive_ram_block ram_block1a21(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "rom";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = 256'h000000000000F361F987E3660220C402408200A0148841042083121125DB1358;

cycloneive_ram_block ram_block1a30(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "rom";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = 256'h000000000001009E007800804331021000000C06C00000061000181980000000;

cycloneive_ram_block ram_block1a29(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "rom";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = 256'h0000000000010098006000005804F0400000000000060016A021C38008404800;

cycloneive_ram_block ram_block1a28(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "rom";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = 256'h0000000000000E9E00780080DCCC324812288E06C0271449B211A4667801C81C;

cycloneive_ram_block ram_block1a27(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "rom";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = 256'h0000000000010000000000001B340240000020048004001090219819B801801C;

cycloneive_ram_block ram_block1a26(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "rom";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = 256'h000000000000002002800508C00441000000101000000000800000000800000A;

cycloneive_ram_block ram_block1a25(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "rom";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = 256'h00000000000003120048089015D810413871C403607438E308586CACC0000000;

cycloneive_ram_block ram_block1a24(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "rom";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = 256'h000000000000030000000890100441001830D000003018638018010018010100;

cycloneive_ram_block ram_block1a23(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "rom";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = 256'h000000000000071204481891C44410012041040360402080984002002800000A;

cycloneive_ram_block ram_block1a22(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "rom";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = 256'h00000000000000000000000011DC0001204110136040208008406EACE801010A;

cycloneive_ram_block ram_block1a20(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "rom";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = 256'h000000000000A37D51F543442222C2200000000A420000041200121124C90118;

cycloneive_ram_block ram_block1a19(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "rom";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = 256'h000000000000F379F9E7E3662220F482408200A0048841042083121125DB5358;

cycloneive_ram_block ram_block1a18(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "rom";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = 256'h000000000000FBFDF9F7E3662222F6A2408200AA468041043283121135DB1B58;

cycloneive_ram_block ram_block1a17(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "rom";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = 256'h000000000000F361F987E3660222C622408200AA568841043282121135DB1B58;

cycloneive_ram_block ram_block1a31(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "niosII_epcs_boot_rom.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "niosII_epcs:epcs|altsyncram:the_boot_copier_rom|altsyncram_0941:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "rom";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = 256'h0000000000000060018003009CCCC0481228A20000271459A031A4664800001C;

endmodule

module niosII_niosII_epcs_sub (
	clk,
	data_to_cpu_5,
	SCLK_reg1,
	SS_n,
	shift_reg_7,
	reset_n,
	saved_grant_0,
	saved_grant_1,
	out_data_buffer_38,
	src_data_38,
	src_data_39,
	src_data_40,
	data_from_cpu,
	mem_used_1,
	wait_latency_counter_1,
	src_valid,
	src_valid1,
	src_data_46,
	out_data_buffer_65,
	p1_wr_strobe,
	src_payload,
	src_data_66,
	data_to_cpu_0,
	data_to_cpu_1,
	data_to_cpu_2,
	data_to_cpu_3,
	data_to_cpu_4,
	data_to_cpu_11,
	data_to_cpu_13,
	data_to_cpu_12,
	data_to_cpu_14,
	data_to_cpu_15,
	data_to_cpu_10,
	data_to_cpu_9,
	data_to_cpu_8,
	data_to_cpu_7,
	data_to_cpu_6,
	irq_reg1,
	src_payload1,
	epcs_data0)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	data_to_cpu_5;
output 	SCLK_reg1;
output 	SS_n;
output 	shift_reg_7;
input 	reset_n;
input 	saved_grant_0;
input 	saved_grant_1;
input 	out_data_buffer_38;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	[15:0] data_from_cpu;
input 	mem_used_1;
input 	wait_latency_counter_1;
input 	src_valid;
input 	src_valid1;
input 	src_data_46;
input 	out_data_buffer_65;
output 	p1_wr_strobe;
input 	src_payload;
input 	src_data_66;
output 	data_to_cpu_0;
output 	data_to_cpu_1;
output 	data_to_cpu_2;
output 	data_to_cpu_3;
output 	data_to_cpu_4;
output 	data_to_cpu_11;
output 	data_to_cpu_13;
output 	data_to_cpu_12;
output 	data_to_cpu_14;
output 	data_to_cpu_15;
output 	data_to_cpu_10;
output 	data_to_cpu_9;
output 	data_to_cpu_8;
output 	data_to_cpu_7;
output 	data_to_cpu_6;
output 	irq_reg1;
input 	src_payload1;
input 	epcs_data0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \p1_data_wr_strobe~0_combout ;
wire \p1_wr_strobe~0_combout ;
wire \p1_wr_strobe~2_combout ;
wire \wr_strobe~q ;
wire \p1_wr_strobe~3_combout ;
wire \p1_data_wr_strobe~combout ;
wire \data_wr_strobe~q ;
wire \tx_holding_primed~0_combout ;
wire \tx_holding_primed~q ;
wire \Add1~0_combout ;
wire \p1_slowcount[0]~1_combout ;
wire \slowcount[0]~q ;
wire \always11~0_combout ;
wire \state[0]~q ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \Equal9~0_combout ;
wire \state~1_combout ;
wire \state[1]~q ;
wire \Add1~3 ;
wire \Add1~4_combout ;
wire \state[2]~q ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \state[3]~q ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \state~0_combout ;
wire \state[4]~q ;
wire \rx_holding_reg[3]~0_combout ;
wire \transmitting~0_combout ;
wire \transmitting~q ;
wire \p1_slowcount[1]~0_combout ;
wire \slowcount[1]~q ;
wire \Equal2~0_combout ;
wire \MISO_reg~0_combout ;
wire \MISO_reg~q ;
wire \write_tx_holding~combout ;
wire \tx_holding_reg[0]~q ;
wire \shift_reg~11_combout ;
wire \write_shift_reg~0_combout ;
wire \shift_reg[2]~12_combout ;
wire \shift_reg[0]~q ;
wire \tx_holding_reg[1]~q ;
wire \shift_reg~10_combout ;
wire \shift_reg[1]~q ;
wire \tx_holding_reg[2]~q ;
wire \shift_reg~9_combout ;
wire \shift_reg[2]~q ;
wire \tx_holding_reg[3]~q ;
wire \shift_reg~8_combout ;
wire \shift_reg[3]~q ;
wire \tx_holding_reg[4]~q ;
wire \shift_reg~7_combout ;
wire \shift_reg[4]~q ;
wire \tx_holding_reg[5]~q ;
wire \shift_reg~6_combout ;
wire \shift_reg[5]~q ;
wire \rx_holding_reg[5]~q ;
wire \slaveselect_wr_strobe~0_combout ;
wire \epcs_slave_select_holding_reg[5]~q ;
wire \control_wr_strobe~combout ;
wire \SSO_reg~q ;
wire \always6~0_combout ;
wire \epcs_slave_select_reg[5]~q ;
wire \p1_data_to_cpu[5]~18_combout ;
wire \data_to_cpu[5]~0_combout ;
wire \endofpacketvalue_wr_strobe~combout ;
wire \endofpacketvalue_reg[5]~q ;
wire \p1_data_to_cpu[5]~19_combout ;
wire \p1_data_to_cpu[5]~39_combout ;
wire \SCLK_reg~0_combout ;
wire \Equal9~1_combout ;
wire \SCLK_reg~1_combout ;
wire \epcs_slave_select_holding_reg[0]~0_combout ;
wire \epcs_slave_select_holding_reg[0]~q ;
wire \epcs_slave_select_reg[0]~q ;
wire \stateZero~q ;
wire \tx_holding_reg[6]~q ;
wire \shift_reg~5_combout ;
wire \shift_reg[6]~q ;
wire \tx_holding_reg[7]~q ;
wire \shift_reg~4_combout ;
wire \endofpacketvalue_reg[0]~q ;
wire \p1_data_to_cpu[0]~2_combout ;
wire \rx_holding_reg[0]~q ;
wire \data_to_cpu[0]~1_combout ;
wire \p1_data_to_cpu[0]~3_combout ;
wire \endofpacketvalue_reg[1]~q ;
wire \epcs_slave_select_holding_reg[1]~q ;
wire \epcs_slave_select_reg[1]~q ;
wire \p1_data_to_cpu[1]~4_combout ;
wire \rx_holding_reg[1]~q ;
wire \p1_data_to_cpu[1]~5_combout ;
wire \endofpacketvalue_reg[2]~q ;
wire \epcs_slave_select_holding_reg[2]~q ;
wire \epcs_slave_select_reg[2]~q ;
wire \p1_data_to_cpu[2]~6_combout ;
wire \rx_holding_reg[2]~q ;
wire \p1_data_to_cpu[2]~7_combout ;
wire \iROE_reg~q ;
wire \data_to_cpu[4]~2_combout ;
wire \epcs_slave_select_holding_reg[3]~q ;
wire \epcs_slave_select_reg[3]~q ;
wire \status_wr_strobe~combout ;
wire \p1_data_rd_strobe~0_combout ;
wire \p1_rd_strobe~0_combout ;
wire \rd_strobe~q ;
wire \p1_data_rd_strobe~combout ;
wire \data_rd_strobe~q ;
wire \RRDY~0_combout ;
wire \RRDY~q ;
wire \ROE~0_combout ;
wire \ROE~q ;
wire \p1_data_to_cpu[3]~8_combout ;
wire \endofpacketvalue_reg[3]~q ;
wire \p1_data_to_cpu[3]~9_combout ;
wire \rx_holding_reg[3]~q ;
wire \p1_data_to_cpu[3]~10_combout ;
wire \iTOE_reg~q ;
wire \epcs_slave_select_holding_reg[4]~q ;
wire \epcs_slave_select_reg[4]~q ;
wire \TRDY~0_combout ;
wire \TOE~0_combout ;
wire \TOE~q ;
wire \p1_data_to_cpu[4]~11_combout ;
wire \endofpacketvalue_reg[4]~q ;
wire \p1_data_to_cpu[4]~12_combout ;
wire \rx_holding_reg[4]~q ;
wire \p1_data_to_cpu[4]~13_combout ;
wire \p1_data_to_cpu[15]~14_combout ;
wire \endofpacketvalue_reg[11]~q ;
wire \epcs_slave_select_holding_reg[11]~q ;
wire \epcs_slave_select_reg[11]~q ;
wire \p1_data_to_cpu[11]~15_combout ;
wire \endofpacketvalue_reg[13]~q ;
wire \epcs_slave_select_holding_reg[13]~q ;
wire \epcs_slave_select_reg[13]~q ;
wire \p1_data_to_cpu[13]~16_combout ;
wire \endofpacketvalue_reg[12]~q ;
wire \epcs_slave_select_holding_reg[12]~q ;
wire \epcs_slave_select_reg[12]~q ;
wire \p1_data_to_cpu[12]~17_combout ;
wire \endofpacketvalue_reg[14]~q ;
wire \epcs_slave_select_holding_reg[14]~q ;
wire \epcs_slave_select_reg[14]~q ;
wire \p1_data_to_cpu[14]~20_combout ;
wire \endofpacketvalue_reg[15]~q ;
wire \epcs_slave_select_holding_reg[15]~q ;
wire \epcs_slave_select_reg[15]~q ;
wire \p1_data_to_cpu[15]~21_combout ;
wire \endofpacketvalue_reg[10]~q ;
wire \epcs_slave_select_holding_reg[10]~q ;
wire \epcs_slave_select_reg[10]~q ;
wire \p1_data_to_cpu[10]~22_combout ;
wire \p1_data_to_cpu[10]~23_combout ;
wire \p1_data_to_cpu[10]~24_combout ;
wire \endofpacketvalue_reg[9]~q ;
wire \epcs_slave_select_holding_reg[9]~q ;
wire \epcs_slave_select_reg[9]~q ;
wire \p1_data_to_cpu[9]~25_combout ;
wire \data_to_cpu[8]~3_combout ;
wire \iEOP_reg~q ;
wire \EOP~0_combout ;
wire \endofpacketvalue_reg[8]~q ;
wire \EOP~1_combout ;
wire \EOP~2_combout ;
wire \EOP~3_combout ;
wire \EOP~4_combout ;
wire \endofpacketvalue_reg[7]~q ;
wire \endofpacketvalue_reg[6]~q ;
wire \rx_holding_reg[6]~q ;
wire \rx_holding_reg[7]~q ;
wire \EOP~5_combout ;
wire \EOP~6_combout ;
wire \EOP~7_combout ;
wire \EOP~8_combout ;
wire \EOP~9_combout ;
wire \EOP~10_combout ;
wire \EOP~11_combout ;
wire \EOP~12_combout ;
wire \EOP~13_combout ;
wire \EOP~14_combout ;
wire \EOP~15_combout ;
wire \EOP~q ;
wire \p1_data_to_cpu[9]~26_combout ;
wire \p1_data_to_cpu[9]~27_combout ;
wire \p1_data_to_cpu[9]~28_combout ;
wire \epcs_slave_select_holding_reg[8]~q ;
wire \epcs_slave_select_reg[8]~q ;
wire \p1_data_to_cpu[8]~29_combout ;
wire \iE_reg~q ;
wire \E~combout ;
wire \p1_data_to_cpu[8]~30_combout ;
wire \p1_data_to_cpu[8]~31_combout ;
wire \p1_data_to_cpu[8]~32_combout ;
wire \iRRDY_reg~q ;
wire \epcs_slave_select_holding_reg[7]~q ;
wire \epcs_slave_select_reg[7]~q ;
wire \p1_data_to_cpu[7]~33_combout ;
wire \p1_data_to_cpu[7]~34_combout ;
wire \p1_data_to_cpu[7]~35_combout ;
wire \iTRDY_reg~q ;
wire \epcs_slave_select_holding_reg[6]~q ;
wire \epcs_slave_select_reg[6]~q ;
wire \p1_data_to_cpu[6]~36_combout ;
wire \p1_data_to_cpu[6]~37_combout ;
wire \p1_data_to_cpu[6]~38_combout ;
wire \irq_reg~0_combout ;
wire \irq_reg~1_combout ;
wire \irq_reg~2_combout ;
wire \irq_reg~3_combout ;


dffeas \data_to_cpu[5] (
	.clk(clk),
	.d(\data_to_cpu[5]~0_combout ),
	.asdata(\p1_data_to_cpu[5]~39_combout ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(src_data_39),
	.ena(vcc),
	.q(data_to_cpu_5),
	.prn(vcc));
defparam \data_to_cpu[5] .is_wysiwyg = "true";
defparam \data_to_cpu[5] .power_up = "low";

dffeas SCLK_reg(
	.clk(clk),
	.d(\SCLK_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(SCLK_reg1),
	.prn(vcc));
defparam SCLK_reg.is_wysiwyg = "true";
defparam SCLK_reg.power_up = "low";

cycloneive_lcell_comb \SS_n~0 (
	.dataa(\epcs_slave_select_reg[0]~q ),
	.datab(\stateZero~q ),
	.datac(\transmitting~q ),
	.datad(\SSO_reg~q ),
	.cin(gnd),
	.combout(SS_n),
	.cout());
defparam \SS_n~0 .lut_mask = 16'hBFFF;
defparam \SS_n~0 .sum_lutc_input = "datac";

dffeas \shift_reg[7] (
	.clk(clk),
	.d(\shift_reg~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg[2]~12_combout ),
	.q(shift_reg_7),
	.prn(vcc));
defparam \shift_reg[7] .is_wysiwyg = "true";
defparam \shift_reg[7] .power_up = "low";

cycloneive_lcell_comb \p1_wr_strobe~1 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_65),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(p1_wr_strobe),
	.cout());
defparam \p1_wr_strobe~1 .lut_mask = 16'hEEEE;
defparam \p1_wr_strobe~1 .sum_lutc_input = "datac";

dffeas \data_to_cpu[0] (
	.clk(clk),
	.d(\p1_data_to_cpu[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_0),
	.prn(vcc));
defparam \data_to_cpu[0] .is_wysiwyg = "true";
defparam \data_to_cpu[0] .power_up = "low";

dffeas \data_to_cpu[1] (
	.clk(clk),
	.d(\p1_data_to_cpu[1]~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_1),
	.prn(vcc));
defparam \data_to_cpu[1] .is_wysiwyg = "true";
defparam \data_to_cpu[1] .power_up = "low";

dffeas \data_to_cpu[2] (
	.clk(clk),
	.d(\p1_data_to_cpu[2]~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_2),
	.prn(vcc));
defparam \data_to_cpu[2] .is_wysiwyg = "true";
defparam \data_to_cpu[2] .power_up = "low";

dffeas \data_to_cpu[3] (
	.clk(clk),
	.d(\p1_data_to_cpu[3]~10_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_3),
	.prn(vcc));
defparam \data_to_cpu[3] .is_wysiwyg = "true";
defparam \data_to_cpu[3] .power_up = "low";

dffeas \data_to_cpu[4] (
	.clk(clk),
	.d(\p1_data_to_cpu[4]~13_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_4),
	.prn(vcc));
defparam \data_to_cpu[4] .is_wysiwyg = "true";
defparam \data_to_cpu[4] .power_up = "low";

dffeas \data_to_cpu[11] (
	.clk(clk),
	.d(\p1_data_to_cpu[11]~15_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_11),
	.prn(vcc));
defparam \data_to_cpu[11] .is_wysiwyg = "true";
defparam \data_to_cpu[11] .power_up = "low";

dffeas \data_to_cpu[13] (
	.clk(clk),
	.d(\p1_data_to_cpu[13]~16_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_13),
	.prn(vcc));
defparam \data_to_cpu[13] .is_wysiwyg = "true";
defparam \data_to_cpu[13] .power_up = "low";

dffeas \data_to_cpu[12] (
	.clk(clk),
	.d(\p1_data_to_cpu[12]~17_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_12),
	.prn(vcc));
defparam \data_to_cpu[12] .is_wysiwyg = "true";
defparam \data_to_cpu[12] .power_up = "low";

dffeas \data_to_cpu[14] (
	.clk(clk),
	.d(\p1_data_to_cpu[14]~20_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_14),
	.prn(vcc));
defparam \data_to_cpu[14] .is_wysiwyg = "true";
defparam \data_to_cpu[14] .power_up = "low";

dffeas \data_to_cpu[15] (
	.clk(clk),
	.d(\p1_data_to_cpu[15]~21_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_15),
	.prn(vcc));
defparam \data_to_cpu[15] .is_wysiwyg = "true";
defparam \data_to_cpu[15] .power_up = "low";

dffeas \data_to_cpu[10] (
	.clk(clk),
	.d(\p1_data_to_cpu[10]~24_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_10),
	.prn(vcc));
defparam \data_to_cpu[10] .is_wysiwyg = "true";
defparam \data_to_cpu[10] .power_up = "low";

dffeas \data_to_cpu[9] (
	.clk(clk),
	.d(\p1_data_to_cpu[9]~28_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_9),
	.prn(vcc));
defparam \data_to_cpu[9] .is_wysiwyg = "true";
defparam \data_to_cpu[9] .power_up = "low";

dffeas \data_to_cpu[8] (
	.clk(clk),
	.d(\p1_data_to_cpu[8]~32_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_8),
	.prn(vcc));
defparam \data_to_cpu[8] .is_wysiwyg = "true";
defparam \data_to_cpu[8] .power_up = "low";

dffeas \data_to_cpu[7] (
	.clk(clk),
	.d(\p1_data_to_cpu[7]~35_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_7),
	.prn(vcc));
defparam \data_to_cpu[7] .is_wysiwyg = "true";
defparam \data_to_cpu[7] .power_up = "low";

dffeas \data_to_cpu[6] (
	.clk(clk),
	.d(\p1_data_to_cpu[6]~38_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_cpu_6),
	.prn(vcc));
defparam \data_to_cpu[6] .is_wysiwyg = "true";
defparam \data_to_cpu[6] .power_up = "low";

dffeas irq_reg(
	.clk(clk),
	.d(\irq_reg~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(irq_reg1),
	.prn(vcc));
defparam irq_reg.is_wysiwyg = "true";
defparam irq_reg.power_up = "low";

cycloneive_lcell_comb \p1_data_wr_strobe~0 (
	.dataa(src_payload),
	.datab(saved_grant_1),
	.datac(out_data_buffer_38),
	.datad(src_data_40),
	.cin(gnd),
	.combout(\p1_data_wr_strobe~0_combout ),
	.cout());
defparam \p1_data_wr_strobe~0 .lut_mask = 16'hFEFF;
defparam \p1_data_wr_strobe~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_wr_strobe~0 (
	.dataa(src_data_46),
	.datab(src_valid),
	.datac(src_valid1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\p1_wr_strobe~0_combout ),
	.cout());
defparam \p1_wr_strobe~0 .lut_mask = 16'hFEFF;
defparam \p1_wr_strobe~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_wr_strobe~2 (
	.dataa(\p1_wr_strobe~0_combout ),
	.datab(p1_wr_strobe),
	.datac(\wr_strobe~q ),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\p1_wr_strobe~2_combout ),
	.cout());
defparam \p1_wr_strobe~2 .lut_mask = 16'hEFFF;
defparam \p1_wr_strobe~2 .sum_lutc_input = "datac";

dffeas wr_strobe(
	.clk(clk),
	.d(\p1_wr_strobe~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_strobe~q ),
	.prn(vcc));
defparam wr_strobe.is_wysiwyg = "true";
defparam wr_strobe.power_up = "low";

cycloneive_lcell_comb \p1_wr_strobe~3 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_65),
	.datac(\wr_strobe~q ),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\p1_wr_strobe~3_combout ),
	.cout());
defparam \p1_wr_strobe~3 .lut_mask = 16'hEFFF;
defparam \p1_wr_strobe~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb p1_data_wr_strobe(
	.dataa(\p1_data_wr_strobe~0_combout ),
	.datab(\p1_wr_strobe~0_combout ),
	.datac(\p1_wr_strobe~3_combout ),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_wr_strobe~combout ),
	.cout());
defparam p1_data_wr_strobe.lut_mask = 16'hFEFF;
defparam p1_data_wr_strobe.sum_lutc_input = "datac";

dffeas data_wr_strobe(
	.clk(clk),
	.d(\p1_data_wr_strobe~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_wr_strobe~q ),
	.prn(vcc));
defparam data_wr_strobe.is_wysiwyg = "true";
defparam data_wr_strobe.power_up = "low";

cycloneive_lcell_comb \tx_holding_primed~0 (
	.dataa(\data_wr_strobe~q ),
	.datab(\transmitting~q ),
	.datac(\tx_holding_primed~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\tx_holding_primed~0_combout ),
	.cout());
defparam \tx_holding_primed~0 .lut_mask = 16'hFEFE;
defparam \tx_holding_primed~0 .sum_lutc_input = "datac";

dffeas tx_holding_primed(
	.clk(clk),
	.d(\tx_holding_primed~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tx_holding_primed~q ),
	.prn(vcc));
defparam tx_holding_primed.is_wysiwyg = "true";
defparam tx_holding_primed.power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(\state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
defparam \Add1~0 .lut_mask = 16'h55AA;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_slowcount[0]~1 (
	.dataa(\transmitting~q ),
	.datab(gnd),
	.datac(\slowcount[1]~q ),
	.datad(\slowcount[0]~q ),
	.cin(gnd),
	.combout(\p1_slowcount[0]~1_combout ),
	.cout());
defparam \p1_slowcount[0]~1 .lut_mask = 16'hAFFF;
defparam \p1_slowcount[0]~1 .sum_lutc_input = "datac";

dffeas \slowcount[0] (
	.clk(clk),
	.d(\p1_slowcount[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\slowcount[0]~q ),
	.prn(vcc));
defparam \slowcount[0] .is_wysiwyg = "true";
defparam \slowcount[0] .power_up = "low";

cycloneive_lcell_comb \always11~0 (
	.dataa(\transmitting~q ),
	.datab(\slowcount[1]~q ),
	.datac(gnd),
	.datad(\slowcount[0]~q ),
	.cin(gnd),
	.combout(\always11~0_combout ),
	.cout());
defparam \always11~0 .lut_mask = 16'hEEFF;
defparam \always11~0 .sum_lutc_input = "datac";

dffeas \state[0] (
	.clk(clk),
	.d(\Add1~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\state[0]~q ),
	.prn(vcc));
defparam \state[0] .is_wysiwyg = "true";
defparam \state[0] .power_up = "low";

cycloneive_lcell_comb \Add1~2 (
	.dataa(\state[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
defparam \Add1~2 .lut_mask = 16'h5A5F;
defparam \Add1~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Equal9~0 (
	.dataa(gnd),
	.datab(\state[3]~q ),
	.datac(\state[2]~q ),
	.datad(\state[1]~q ),
	.cin(gnd),
	.combout(\Equal9~0_combout ),
	.cout());
defparam \Equal9~0 .lut_mask = 16'h3FFF;
defparam \Equal9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~1 (
	.dataa(\Add1~2_combout ),
	.datab(\state[0]~q ),
	.datac(\state[4]~q ),
	.datad(\Equal9~0_combout ),
	.cin(gnd),
	.combout(\state~1_combout ),
	.cout());
defparam \state~1 .lut_mask = 16'hBFFF;
defparam \state~1 .sum_lutc_input = "datac";

dffeas \state[1] (
	.clk(clk),
	.d(\state~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\state[1]~q ),
	.prn(vcc));
defparam \state[1] .is_wysiwyg = "true";
defparam \state[1] .power_up = "low";

cycloneive_lcell_comb \Add1~4 (
	.dataa(\state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
defparam \Add1~4 .lut_mask = 16'h5AAF;
defparam \Add1~4 .sum_lutc_input = "cin";

dffeas \state[2] (
	.clk(clk),
	.d(\Add1~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\state[2]~q ),
	.prn(vcc));
defparam \state[2] .is_wysiwyg = "true";
defparam \state[2] .power_up = "low";

cycloneive_lcell_comb \Add1~6 (
	.dataa(\state[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";

dffeas \state[3] (
	.clk(clk),
	.d(\Add1~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\state[3]~q ),
	.prn(vcc));
defparam \state[3] .is_wysiwyg = "true";
defparam \state[3] .power_up = "low";

cycloneive_lcell_comb \Add1~8 (
	.dataa(\state[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout());
defparam \Add1~8 .lut_mask = 16'h5A5A;
defparam \Add1~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \state~0 (
	.dataa(\Add1~8_combout ),
	.datab(\state[0]~q ),
	.datac(\state[4]~q ),
	.datad(\Equal9~0_combout ),
	.cin(gnd),
	.combout(\state~0_combout ),
	.cout());
defparam \state~0 .lut_mask = 16'hBFFF;
defparam \state~0 .sum_lutc_input = "datac";

dffeas \state[4] (
	.clk(clk),
	.d(\state~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\state[4]~q ),
	.prn(vcc));
defparam \state[4] .is_wysiwyg = "true";
defparam \state[4] .power_up = "low";

cycloneive_lcell_comb \rx_holding_reg[3]~0 (
	.dataa(\Equal2~0_combout ),
	.datab(\state[0]~q ),
	.datac(\state[4]~q ),
	.datad(\Equal9~0_combout ),
	.cin(gnd),
	.combout(\rx_holding_reg[3]~0_combout ),
	.cout());
defparam \rx_holding_reg[3]~0 .lut_mask = 16'hFFFE;
defparam \rx_holding_reg[3]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \transmitting~0 (
	.dataa(\transmitting~q ),
	.datab(\tx_holding_primed~q ),
	.datac(gnd),
	.datad(\rx_holding_reg[3]~0_combout ),
	.cin(gnd),
	.combout(\transmitting~0_combout ),
	.cout());
defparam \transmitting~0 .lut_mask = 16'hEEFF;
defparam \transmitting~0 .sum_lutc_input = "datac";

dffeas transmitting(
	.clk(clk),
	.d(\transmitting~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\transmitting~q ),
	.prn(vcc));
defparam transmitting.is_wysiwyg = "true";
defparam transmitting.power_up = "low";

cycloneive_lcell_comb \p1_slowcount[1]~0 (
	.dataa(\transmitting~q ),
	.datab(\slowcount[0]~q ),
	.datac(gnd),
	.datad(\slowcount[1]~q ),
	.cin(gnd),
	.combout(\p1_slowcount[1]~0_combout ),
	.cout());
defparam \p1_slowcount[1]~0 .lut_mask = 16'hEEFF;
defparam \p1_slowcount[1]~0 .sum_lutc_input = "datac";

dffeas \slowcount[1] (
	.clk(clk),
	.d(\p1_slowcount[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\slowcount[1]~q ),
	.prn(vcc));
defparam \slowcount[1] .is_wysiwyg = "true";
defparam \slowcount[1] .power_up = "low";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(\slowcount[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\slowcount[0]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hAAFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MISO_reg~0 (
	.dataa(\MISO_reg~q ),
	.datab(epcs_data0),
	.datac(\Equal2~0_combout ),
	.datad(SCLK_reg1),
	.cin(gnd),
	.combout(\MISO_reg~0_combout ),
	.cout());
defparam \MISO_reg~0 .lut_mask = 16'hEFFE;
defparam \MISO_reg~0 .sum_lutc_input = "datac";

dffeas MISO_reg(
	.clk(clk),
	.d(\MISO_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\MISO_reg~q ),
	.prn(vcc));
defparam MISO_reg.is_wysiwyg = "true";
defparam MISO_reg.power_up = "low";

cycloneive_lcell_comb write_tx_holding(
	.dataa(\data_wr_strobe~q ),
	.datab(gnd),
	.datac(\transmitting~q ),
	.datad(\tx_holding_primed~q ),
	.cin(gnd),
	.combout(\write_tx_holding~combout ),
	.cout());
defparam write_tx_holding.lut_mask = 16'hAFFF;
defparam write_tx_holding.sum_lutc_input = "datac";

dffeas \tx_holding_reg[0] (
	.clk(clk),
	.d(data_from_cpu[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_tx_holding~combout ),
	.q(\tx_holding_reg[0]~q ),
	.prn(vcc));
defparam \tx_holding_reg[0] .is_wysiwyg = "true";
defparam \tx_holding_reg[0] .power_up = "low";

cycloneive_lcell_comb \shift_reg~11 (
	.dataa(\MISO_reg~q ),
	.datab(\tx_holding_reg[0]~q ),
	.datac(SCLK_reg1),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\shift_reg~11_combout ),
	.cout());
defparam \shift_reg~11 .lut_mask = 16'hEFFE;
defparam \shift_reg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_shift_reg~0 (
	.dataa(\tx_holding_primed~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\transmitting~q ),
	.cin(gnd),
	.combout(\write_shift_reg~0_combout ),
	.cout());
defparam \write_shift_reg~0 .lut_mask = 16'hAAFF;
defparam \write_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shift_reg[2]~12 (
	.dataa(\slowcount[1]~q ),
	.datab(\slowcount[0]~q ),
	.datac(SCLK_reg1),
	.datad(\write_shift_reg~0_combout ),
	.cin(gnd),
	.combout(\shift_reg[2]~12_combout ),
	.cout());
defparam \shift_reg[2]~12 .lut_mask = 16'hFFFB;
defparam \shift_reg[2]~12 .sum_lutc_input = "datac";

dffeas \shift_reg[0] (
	.clk(clk),
	.d(\shift_reg~11_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg[2]~12_combout ),
	.q(\shift_reg[0]~q ),
	.prn(vcc));
defparam \shift_reg[0] .is_wysiwyg = "true";
defparam \shift_reg[0] .power_up = "low";

dffeas \tx_holding_reg[1] (
	.clk(clk),
	.d(data_from_cpu[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_tx_holding~combout ),
	.q(\tx_holding_reg[1]~q ),
	.prn(vcc));
defparam \tx_holding_reg[1] .is_wysiwyg = "true";
defparam \tx_holding_reg[1] .power_up = "low";

cycloneive_lcell_comb \shift_reg~10 (
	.dataa(\shift_reg[0]~q ),
	.datab(\tx_holding_reg[1]~q ),
	.datac(SCLK_reg1),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\shift_reg~10_combout ),
	.cout());
defparam \shift_reg~10 .lut_mask = 16'hEFFE;
defparam \shift_reg~10 .sum_lutc_input = "datac";

dffeas \shift_reg[1] (
	.clk(clk),
	.d(\shift_reg~10_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg[2]~12_combout ),
	.q(\shift_reg[1]~q ),
	.prn(vcc));
defparam \shift_reg[1] .is_wysiwyg = "true";
defparam \shift_reg[1] .power_up = "low";

dffeas \tx_holding_reg[2] (
	.clk(clk),
	.d(data_from_cpu[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_tx_holding~combout ),
	.q(\tx_holding_reg[2]~q ),
	.prn(vcc));
defparam \tx_holding_reg[2] .is_wysiwyg = "true";
defparam \tx_holding_reg[2] .power_up = "low";

cycloneive_lcell_comb \shift_reg~9 (
	.dataa(\shift_reg[1]~q ),
	.datab(\tx_holding_reg[2]~q ),
	.datac(SCLK_reg1),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\shift_reg~9_combout ),
	.cout());
defparam \shift_reg~9 .lut_mask = 16'hEFFE;
defparam \shift_reg~9 .sum_lutc_input = "datac";

dffeas \shift_reg[2] (
	.clk(clk),
	.d(\shift_reg~9_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg[2]~12_combout ),
	.q(\shift_reg[2]~q ),
	.prn(vcc));
defparam \shift_reg[2] .is_wysiwyg = "true";
defparam \shift_reg[2] .power_up = "low";

dffeas \tx_holding_reg[3] (
	.clk(clk),
	.d(data_from_cpu[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_tx_holding~combout ),
	.q(\tx_holding_reg[3]~q ),
	.prn(vcc));
defparam \tx_holding_reg[3] .is_wysiwyg = "true";
defparam \tx_holding_reg[3] .power_up = "low";

cycloneive_lcell_comb \shift_reg~8 (
	.dataa(\shift_reg[2]~q ),
	.datab(\tx_holding_reg[3]~q ),
	.datac(SCLK_reg1),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\shift_reg~8_combout ),
	.cout());
defparam \shift_reg~8 .lut_mask = 16'hEFFE;
defparam \shift_reg~8 .sum_lutc_input = "datac";

dffeas \shift_reg[3] (
	.clk(clk),
	.d(\shift_reg~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg[2]~12_combout ),
	.q(\shift_reg[3]~q ),
	.prn(vcc));
defparam \shift_reg[3] .is_wysiwyg = "true";
defparam \shift_reg[3] .power_up = "low";

dffeas \tx_holding_reg[4] (
	.clk(clk),
	.d(data_from_cpu[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_tx_holding~combout ),
	.q(\tx_holding_reg[4]~q ),
	.prn(vcc));
defparam \tx_holding_reg[4] .is_wysiwyg = "true";
defparam \tx_holding_reg[4] .power_up = "low";

cycloneive_lcell_comb \shift_reg~7 (
	.dataa(\shift_reg[3]~q ),
	.datab(\tx_holding_reg[4]~q ),
	.datac(SCLK_reg1),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\shift_reg~7_combout ),
	.cout());
defparam \shift_reg~7 .lut_mask = 16'hEFFE;
defparam \shift_reg~7 .sum_lutc_input = "datac";

dffeas \shift_reg[4] (
	.clk(clk),
	.d(\shift_reg~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg[2]~12_combout ),
	.q(\shift_reg[4]~q ),
	.prn(vcc));
defparam \shift_reg[4] .is_wysiwyg = "true";
defparam \shift_reg[4] .power_up = "low";

dffeas \tx_holding_reg[5] (
	.clk(clk),
	.d(data_from_cpu[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_tx_holding~combout ),
	.q(\tx_holding_reg[5]~q ),
	.prn(vcc));
defparam \tx_holding_reg[5] .is_wysiwyg = "true";
defparam \tx_holding_reg[5] .power_up = "low";

cycloneive_lcell_comb \shift_reg~6 (
	.dataa(\shift_reg[4]~q ),
	.datab(\tx_holding_reg[5]~q ),
	.datac(SCLK_reg1),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\shift_reg~6_combout ),
	.cout());
defparam \shift_reg~6 .lut_mask = 16'hEFFE;
defparam \shift_reg~6 .sum_lutc_input = "datac";

dffeas \shift_reg[5] (
	.clk(clk),
	.d(\shift_reg~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg[2]~12_combout ),
	.q(\shift_reg[5]~q ),
	.prn(vcc));
defparam \shift_reg[5] .is_wysiwyg = "true";
defparam \shift_reg[5] .power_up = "low";

dffeas \rx_holding_reg[5] (
	.clk(clk),
	.d(\shift_reg[5]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_holding_reg[3]~0_combout ),
	.q(\rx_holding_reg[5]~q ),
	.prn(vcc));
defparam \rx_holding_reg[5] .is_wysiwyg = "true";
defparam \rx_holding_reg[5] .power_up = "low";

cycloneive_lcell_comb \slaveselect_wr_strobe~0 (
	.dataa(src_data_38),
	.datab(src_data_40),
	.datac(\wr_strobe~q ),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\slaveselect_wr_strobe~0_combout ),
	.cout());
defparam \slaveselect_wr_strobe~0 .lut_mask = 16'hFEFF;
defparam \slaveselect_wr_strobe~0 .sum_lutc_input = "datac";

dffeas \epcs_slave_select_holding_reg[5] (
	.clk(clk),
	.d(data_from_cpu[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[5]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[5] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[5] .power_up = "low";

cycloneive_lcell_comb control_wr_strobe(
	.dataa(src_data_38),
	.datab(\wr_strobe~q ),
	.datac(src_data_39),
	.datad(src_data_40),
	.cin(gnd),
	.combout(\control_wr_strobe~combout ),
	.cout());
defparam control_wr_strobe.lut_mask = 16'hFEFF;
defparam control_wr_strobe.sum_lutc_input = "datac";

dffeas SSO_reg(
	.clk(clk),
	.d(data_from_cpu[10]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\SSO_reg~q ),
	.prn(vcc));
defparam SSO_reg.is_wysiwyg = "true";
defparam SSO_reg.power_up = "low";

cycloneive_lcell_comb \always6~0 (
	.dataa(\write_shift_reg~0_combout ),
	.datab(\control_wr_strobe~combout ),
	.datac(data_from_cpu[10]),
	.datad(\SSO_reg~q ),
	.cin(gnd),
	.combout(\always6~0_combout ),
	.cout());
defparam \always6~0 .lut_mask = 16'hFEFF;
defparam \always6~0 .sum_lutc_input = "datac";

dffeas \epcs_slave_select_reg[5] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[5]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[5]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[5] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[5] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[5]~18 (
	.dataa(src_data_38),
	.datab(src_data_40),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p1_data_to_cpu[5]~18_combout ),
	.cout());
defparam \p1_data_to_cpu[5]~18 .lut_mask = 16'hEEEE;
defparam \p1_data_to_cpu[5]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_to_cpu[5]~0 (
	.dataa(\rx_holding_reg[5]~q ),
	.datab(\epcs_slave_select_reg[5]~q ),
	.datac(gnd),
	.datad(\p1_data_to_cpu[5]~18_combout ),
	.cin(gnd),
	.combout(\data_to_cpu[5]~0_combout ),
	.cout());
defparam \data_to_cpu[5]~0 .lut_mask = 16'hAACC;
defparam \data_to_cpu[5]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb endofpacketvalue_wr_strobe(
	.dataa(src_data_40),
	.datab(\wr_strobe~q ),
	.datac(src_data_39),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\endofpacketvalue_wr_strobe~combout ),
	.cout());
defparam endofpacketvalue_wr_strobe.lut_mask = 16'hFEFF;
defparam endofpacketvalue_wr_strobe.sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[5] (
	.clk(clk),
	.d(data_from_cpu[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[5]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[5] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[5] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[5]~19 (
	.dataa(\endofpacketvalue_reg[5]~q ),
	.datab(src_data_40),
	.datac(\transmitting~q ),
	.datad(\tx_holding_primed~q ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[5]~19_combout ),
	.cout());
defparam \p1_data_to_cpu[5]~19 .lut_mask = 16'h8BFF;
defparam \p1_data_to_cpu[5]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[5]~39 (
	.dataa(src_data_38),
	.datab(src_data_40),
	.datac(\rx_holding_reg[5]~q ),
	.datad(\p1_data_to_cpu[5]~19_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[5]~39_combout ),
	.cout());
defparam \p1_data_to_cpu[5]~39 .lut_mask = 16'hFFD8;
defparam \p1_data_to_cpu[5]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \SCLK_reg~0 (
	.dataa(\transmitting~q ),
	.datab(\state[0]~q ),
	.datac(\state[4]~q ),
	.datad(\Equal9~0_combout ),
	.cin(gnd),
	.combout(\SCLK_reg~0_combout ),
	.cout());
defparam \SCLK_reg~0 .lut_mask = 16'hFEFF;
defparam \SCLK_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal9~1 (
	.dataa(\state[0]~q ),
	.datab(\state[4]~q ),
	.datac(\Equal9~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal9~1_combout ),
	.cout());
defparam \Equal9~1 .lut_mask = 16'h7F7F;
defparam \Equal9~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \SCLK_reg~1 (
	.dataa(SCLK_reg1),
	.datab(\SCLK_reg~0_combout ),
	.datac(\Equal9~1_combout ),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\SCLK_reg~1_combout ),
	.cout());
defparam \SCLK_reg~1 .lut_mask = 16'hF9F6;
defparam \SCLK_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \epcs_slave_select_holding_reg[0]~0 (
	.dataa(data_from_cpu[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\epcs_slave_select_holding_reg[0]~0_combout ),
	.cout());
defparam \epcs_slave_select_holding_reg[0]~0 .lut_mask = 16'h5555;
defparam \epcs_slave_select_holding_reg[0]~0 .sum_lutc_input = "datac";

dffeas \epcs_slave_select_holding_reg[0] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[0]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[0] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[0] .power_up = "low";

dffeas \epcs_slave_select_reg[0] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[0]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[0] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[0] .power_up = "low";

dffeas stateZero(
	.clk(clk),
	.d(\Equal9~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always11~0_combout ),
	.q(\stateZero~q ),
	.prn(vcc));
defparam stateZero.is_wysiwyg = "true";
defparam stateZero.power_up = "low";

dffeas \tx_holding_reg[6] (
	.clk(clk),
	.d(data_from_cpu[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_tx_holding~combout ),
	.q(\tx_holding_reg[6]~q ),
	.prn(vcc));
defparam \tx_holding_reg[6] .is_wysiwyg = "true";
defparam \tx_holding_reg[6] .power_up = "low";

cycloneive_lcell_comb \shift_reg~5 (
	.dataa(\shift_reg[5]~q ),
	.datab(\tx_holding_reg[6]~q ),
	.datac(SCLK_reg1),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\shift_reg~5_combout ),
	.cout());
defparam \shift_reg~5 .lut_mask = 16'hEFFE;
defparam \shift_reg~5 .sum_lutc_input = "datac";

dffeas \shift_reg[6] (
	.clk(clk),
	.d(\shift_reg~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg[2]~12_combout ),
	.q(\shift_reg[6]~q ),
	.prn(vcc));
defparam \shift_reg[6] .is_wysiwyg = "true";
defparam \shift_reg[6] .power_up = "low";

dffeas \tx_holding_reg[7] (
	.clk(clk),
	.d(data_from_cpu[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_tx_holding~combout ),
	.q(\tx_holding_reg[7]~q ),
	.prn(vcc));
defparam \tx_holding_reg[7] .is_wysiwyg = "true";
defparam \tx_holding_reg[7] .power_up = "low";

cycloneive_lcell_comb \shift_reg~4 (
	.dataa(\shift_reg[6]~q ),
	.datab(\tx_holding_reg[7]~q ),
	.datac(SCLK_reg1),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\shift_reg~4_combout ),
	.cout());
defparam \shift_reg~4 .lut_mask = 16'hEFFE;
defparam \shift_reg~4 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[0] (
	.clk(clk),
	.d(data_from_cpu[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[0]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[0] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[0] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[0]~2 (
	.dataa(\endofpacketvalue_reg[0]~q ),
	.datab(src_data_39),
	.datac(gnd),
	.datad(\epcs_slave_select_reg[0]~q ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[0]~2_combout ),
	.cout());
defparam \p1_data_to_cpu[0]~2 .lut_mask = 16'h88BB;
defparam \p1_data_to_cpu[0]~2 .sum_lutc_input = "datac";

dffeas \rx_holding_reg[0] (
	.clk(clk),
	.d(\shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_holding_reg[3]~0_combout ),
	.q(\rx_holding_reg[0]~q ),
	.prn(vcc));
defparam \rx_holding_reg[0] .is_wysiwyg = "true";
defparam \rx_holding_reg[0] .power_up = "low";

cycloneive_lcell_comb \data_to_cpu[0]~1 (
	.dataa(gnd),
	.datab(src_data_39),
	.datac(src_data_38),
	.datad(src_data_40),
	.cin(gnd),
	.combout(\data_to_cpu[0]~1_combout ),
	.cout());
defparam \data_to_cpu[0]~1 .lut_mask = 16'hC33C;
defparam \data_to_cpu[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[0]~3 (
	.dataa(src_data_40),
	.datab(\p1_data_to_cpu[0]~2_combout ),
	.datac(\rx_holding_reg[0]~q ),
	.datad(\data_to_cpu[0]~1_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[0]~3_combout ),
	.cout());
defparam \p1_data_to_cpu[0]~3 .lut_mask = 16'hFAFC;
defparam \p1_data_to_cpu[0]~3 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[1] (
	.clk(clk),
	.d(data_from_cpu[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[1]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[1] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[1] .power_up = "low";

dffeas \epcs_slave_select_holding_reg[1] (
	.clk(clk),
	.d(data_from_cpu[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[1]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[1] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[1] .power_up = "low";

dffeas \epcs_slave_select_reg[1] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[1]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[1]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[1] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[1] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[1]~4 (
	.dataa(\endofpacketvalue_reg[1]~q ),
	.datab(\epcs_slave_select_reg[1]~q ),
	.datac(gnd),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[1]~4_combout ),
	.cout());
defparam \p1_data_to_cpu[1]~4 .lut_mask = 16'hAACC;
defparam \p1_data_to_cpu[1]~4 .sum_lutc_input = "datac";

dffeas \rx_holding_reg[1] (
	.clk(clk),
	.d(\shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_holding_reg[3]~0_combout ),
	.q(\rx_holding_reg[1]~q ),
	.prn(vcc));
defparam \rx_holding_reg[1] .is_wysiwyg = "true";
defparam \rx_holding_reg[1] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[1]~5 (
	.dataa(src_data_40),
	.datab(\p1_data_to_cpu[1]~4_combout ),
	.datac(\rx_holding_reg[1]~q ),
	.datad(\data_to_cpu[0]~1_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[1]~5_combout ),
	.cout());
defparam \p1_data_to_cpu[1]~5 .lut_mask = 16'hFAFC;
defparam \p1_data_to_cpu[1]~5 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[2] (
	.clk(clk),
	.d(data_from_cpu[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[2]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[2] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[2] .power_up = "low";

dffeas \epcs_slave_select_holding_reg[2] (
	.clk(clk),
	.d(data_from_cpu[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[2]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[2] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[2] .power_up = "low";

dffeas \epcs_slave_select_reg[2] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[2]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[2]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[2] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[2] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[2]~6 (
	.dataa(\endofpacketvalue_reg[2]~q ),
	.datab(\epcs_slave_select_reg[2]~q ),
	.datac(gnd),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[2]~6_combout ),
	.cout());
defparam \p1_data_to_cpu[2]~6 .lut_mask = 16'hAACC;
defparam \p1_data_to_cpu[2]~6 .sum_lutc_input = "datac";

dffeas \rx_holding_reg[2] (
	.clk(clk),
	.d(\shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_holding_reg[3]~0_combout ),
	.q(\rx_holding_reg[2]~q ),
	.prn(vcc));
defparam \rx_holding_reg[2] .is_wysiwyg = "true";
defparam \rx_holding_reg[2] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[2]~7 (
	.dataa(src_data_40),
	.datab(\p1_data_to_cpu[2]~6_combout ),
	.datac(\rx_holding_reg[2]~q ),
	.datad(\data_to_cpu[0]~1_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[2]~7_combout ),
	.cout());
defparam \p1_data_to_cpu[2]~7 .lut_mask = 16'hFAFC;
defparam \p1_data_to_cpu[2]~7 .sum_lutc_input = "datac";

dffeas iROE_reg(
	.clk(clk),
	.d(data_from_cpu[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\iROE_reg~q ),
	.prn(vcc));
defparam iROE_reg.is_wysiwyg = "true";
defparam iROE_reg.power_up = "low";

cycloneive_lcell_comb \data_to_cpu[4]~2 (
	.dataa(src_data_39),
	.datab(src_payload),
	.datac(src_payload1),
	.datad(src_data_40),
	.cin(gnd),
	.combout(\data_to_cpu[4]~2_combout ),
	.cout());
defparam \data_to_cpu[4]~2 .lut_mask = 16'hFAFC;
defparam \data_to_cpu[4]~2 .sum_lutc_input = "datac";

dffeas \epcs_slave_select_holding_reg[3] (
	.clk(clk),
	.d(data_from_cpu[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[3]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[3] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[3] .power_up = "low";

dffeas \epcs_slave_select_reg[3] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[3]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[3]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[3] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[3] .power_up = "low";

cycloneive_lcell_comb status_wr_strobe(
	.dataa(\wr_strobe~q ),
	.datab(src_data_39),
	.datac(src_data_38),
	.datad(src_data_40),
	.cin(gnd),
	.combout(\status_wr_strobe~combout ),
	.cout());
defparam status_wr_strobe.lut_mask = 16'hEFFF;
defparam status_wr_strobe.sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_rd_strobe~0 (
	.dataa(src_payload),
	.datab(src_payload1),
	.datac(src_data_40),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_rd_strobe~0_combout ),
	.cout());
defparam \p1_data_rd_strobe~0 .lut_mask = 16'h7FFF;
defparam \p1_data_rd_strobe~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_rd_strobe~0 (
	.dataa(\p1_wr_strobe~0_combout ),
	.datab(src_data_66),
	.datac(gnd),
	.datad(\rd_strobe~q ),
	.cin(gnd),
	.combout(\p1_rd_strobe~0_combout ),
	.cout());
defparam \p1_rd_strobe~0 .lut_mask = 16'hEEFF;
defparam \p1_rd_strobe~0 .sum_lutc_input = "datac";

dffeas rd_strobe(
	.clk(clk),
	.d(\p1_rd_strobe~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_strobe~q ),
	.prn(vcc));
defparam rd_strobe.is_wysiwyg = "true";
defparam rd_strobe.power_up = "low";

cycloneive_lcell_comb p1_data_rd_strobe(
	.dataa(\p1_wr_strobe~0_combout ),
	.datab(src_data_66),
	.datac(\p1_data_rd_strobe~0_combout ),
	.datad(\rd_strobe~q ),
	.cin(gnd),
	.combout(\p1_data_rd_strobe~combout ),
	.cout());
defparam p1_data_rd_strobe.lut_mask = 16'hFEFF;
defparam p1_data_rd_strobe.sum_lutc_input = "datac";

dffeas data_rd_strobe(
	.clk(clk),
	.d(\p1_data_rd_strobe~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_rd_strobe~q ),
	.prn(vcc));
defparam data_rd_strobe.is_wysiwyg = "true";
defparam data_rd_strobe.power_up = "low";

cycloneive_lcell_comb \RRDY~0 (
	.dataa(\rx_holding_reg[3]~0_combout ),
	.datab(\RRDY~q ),
	.datac(\status_wr_strobe~combout ),
	.datad(\data_rd_strobe~q ),
	.cin(gnd),
	.combout(\RRDY~0_combout ),
	.cout());
defparam \RRDY~0 .lut_mask = 16'hEFFF;
defparam \RRDY~0 .sum_lutc_input = "datac";

dffeas RRDY(
	.clk(clk),
	.d(\RRDY~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\RRDY~q ),
	.prn(vcc));
defparam RRDY.is_wysiwyg = "true";
defparam RRDY.power_up = "low";

cycloneive_lcell_comb \ROE~0 (
	.dataa(\rx_holding_reg[3]~0_combout ),
	.datab(\RRDY~q ),
	.datac(\ROE~q ),
	.datad(\status_wr_strobe~combout ),
	.cin(gnd),
	.combout(\ROE~0_combout ),
	.cout());
defparam \ROE~0 .lut_mask = 16'hFEFF;
defparam \ROE~0 .sum_lutc_input = "datac";

dffeas ROE(
	.clk(clk),
	.d(\ROE~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ROE~q ),
	.prn(vcc));
defparam ROE.is_wysiwyg = "true";
defparam ROE.power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[3]~8 (
	.dataa(\data_to_cpu[4]~2_combout ),
	.datab(\epcs_slave_select_reg[3]~q ),
	.datac(src_data_40),
	.datad(\ROE~q ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[3]~8_combout ),
	.cout());
defparam \p1_data_to_cpu[3]~8 .lut_mask = 16'hFFDE;
defparam \p1_data_to_cpu[3]~8 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[3] (
	.clk(clk),
	.d(data_from_cpu[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[3]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[3] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[3] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[3]~9 (
	.dataa(\iROE_reg~q ),
	.datab(\data_to_cpu[4]~2_combout ),
	.datac(\p1_data_to_cpu[3]~8_combout ),
	.datad(\endofpacketvalue_reg[3]~q ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[3]~9_combout ),
	.cout());
defparam \p1_data_to_cpu[3]~9 .lut_mask = 16'hFFBE;
defparam \p1_data_to_cpu[3]~9 .sum_lutc_input = "datac";

dffeas \rx_holding_reg[3] (
	.clk(clk),
	.d(\shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_holding_reg[3]~0_combout ),
	.q(\rx_holding_reg[3]~q ),
	.prn(vcc));
defparam \rx_holding_reg[3] .is_wysiwyg = "true";
defparam \rx_holding_reg[3] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[3]~10 (
	.dataa(\p1_data_to_cpu[3]~9_combout ),
	.datab(\rx_holding_reg[3]~q ),
	.datac(gnd),
	.datad(\data_to_cpu[0]~1_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[3]~10_combout ),
	.cout());
defparam \p1_data_to_cpu[3]~10 .lut_mask = 16'hAACC;
defparam \p1_data_to_cpu[3]~10 .sum_lutc_input = "datac";

dffeas iTOE_reg(
	.clk(clk),
	.d(data_from_cpu[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\iTOE_reg~q ),
	.prn(vcc));
defparam iTOE_reg.is_wysiwyg = "true";
defparam iTOE_reg.power_up = "low";

dffeas \epcs_slave_select_holding_reg[4] (
	.clk(clk),
	.d(data_from_cpu[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[4]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[4] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[4] .power_up = "low";

dffeas \epcs_slave_select_reg[4] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[4]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[4]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[4] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[4] .power_up = "low";

cycloneive_lcell_comb \TRDY~0 (
	.dataa(\transmitting~q ),
	.datab(\tx_holding_primed~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\TRDY~0_combout ),
	.cout());
defparam \TRDY~0 .lut_mask = 16'hEEEE;
defparam \TRDY~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \TOE~0 (
	.dataa(\TOE~q ),
	.datab(\TRDY~0_combout ),
	.datac(\data_wr_strobe~q ),
	.datad(\status_wr_strobe~combout ),
	.cin(gnd),
	.combout(\TOE~0_combout ),
	.cout());
defparam \TOE~0 .lut_mask = 16'hFEFF;
defparam \TOE~0 .sum_lutc_input = "datac";

dffeas TOE(
	.clk(clk),
	.d(\TOE~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\TOE~q ),
	.prn(vcc));
defparam TOE.is_wysiwyg = "true";
defparam TOE.power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[4]~11 (
	.dataa(\data_to_cpu[4]~2_combout ),
	.datab(\epcs_slave_select_reg[4]~q ),
	.datac(src_data_40),
	.datad(\TOE~q ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[4]~11_combout ),
	.cout());
defparam \p1_data_to_cpu[4]~11 .lut_mask = 16'hFFDE;
defparam \p1_data_to_cpu[4]~11 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[4] (
	.clk(clk),
	.d(data_from_cpu[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[4]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[4] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[4] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[4]~12 (
	.dataa(\iTOE_reg~q ),
	.datab(\data_to_cpu[4]~2_combout ),
	.datac(\p1_data_to_cpu[4]~11_combout ),
	.datad(\endofpacketvalue_reg[4]~q ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[4]~12_combout ),
	.cout());
defparam \p1_data_to_cpu[4]~12 .lut_mask = 16'hFFBE;
defparam \p1_data_to_cpu[4]~12 .sum_lutc_input = "datac";

dffeas \rx_holding_reg[4] (
	.clk(clk),
	.d(\shift_reg[4]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_holding_reg[3]~0_combout ),
	.q(\rx_holding_reg[4]~q ),
	.prn(vcc));
defparam \rx_holding_reg[4] .is_wysiwyg = "true";
defparam \rx_holding_reg[4] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[4]~13 (
	.dataa(\p1_data_to_cpu[4]~12_combout ),
	.datab(\rx_holding_reg[4]~q ),
	.datac(gnd),
	.datad(\data_to_cpu[0]~1_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[4]~13_combout ),
	.cout());
defparam \p1_data_to_cpu[4]~13 .lut_mask = 16'hAACC;
defparam \p1_data_to_cpu[4]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[15]~14 (
	.dataa(src_data_40),
	.datab(gnd),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[15]~14_combout ),
	.cout());
defparam \p1_data_to_cpu[15]~14 .lut_mask = 16'hAFFA;
defparam \p1_data_to_cpu[15]~14 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[11] (
	.clk(clk),
	.d(data_from_cpu[11]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[11]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[11] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[11] .power_up = "low";

dffeas \epcs_slave_select_holding_reg[11] (
	.clk(clk),
	.d(data_from_cpu[11]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[11]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[11] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[11] .power_up = "low";

dffeas \epcs_slave_select_reg[11] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[11]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[11]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[11] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[11] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[11]~15 (
	.dataa(\p1_data_to_cpu[15]~14_combout ),
	.datab(\endofpacketvalue_reg[11]~q ),
	.datac(\epcs_slave_select_reg[11]~q ),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[11]~15_combout ),
	.cout());
defparam \p1_data_to_cpu[11]~15 .lut_mask = 16'hFAFC;
defparam \p1_data_to_cpu[11]~15 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[13] (
	.clk(clk),
	.d(data_from_cpu[13]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[13]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[13] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[13] .power_up = "low";

dffeas \epcs_slave_select_holding_reg[13] (
	.clk(clk),
	.d(data_from_cpu[13]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[13]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[13] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[13] .power_up = "low";

dffeas \epcs_slave_select_reg[13] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[13]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[13]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[13] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[13] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[13]~16 (
	.dataa(\p1_data_to_cpu[15]~14_combout ),
	.datab(\endofpacketvalue_reg[13]~q ),
	.datac(\epcs_slave_select_reg[13]~q ),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[13]~16_combout ),
	.cout());
defparam \p1_data_to_cpu[13]~16 .lut_mask = 16'hFAFC;
defparam \p1_data_to_cpu[13]~16 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[12] (
	.clk(clk),
	.d(data_from_cpu[12]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[12]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[12] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[12] .power_up = "low";

dffeas \epcs_slave_select_holding_reg[12] (
	.clk(clk),
	.d(data_from_cpu[12]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[12]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[12] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[12] .power_up = "low";

dffeas \epcs_slave_select_reg[12] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[12]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[12]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[12] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[12] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[12]~17 (
	.dataa(\p1_data_to_cpu[15]~14_combout ),
	.datab(\endofpacketvalue_reg[12]~q ),
	.datac(\epcs_slave_select_reg[12]~q ),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[12]~17_combout ),
	.cout());
defparam \p1_data_to_cpu[12]~17 .lut_mask = 16'hFAFC;
defparam \p1_data_to_cpu[12]~17 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[14] (
	.clk(clk),
	.d(data_from_cpu[14]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[14]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[14] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[14] .power_up = "low";

dffeas \epcs_slave_select_holding_reg[14] (
	.clk(clk),
	.d(data_from_cpu[14]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[14]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[14] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[14] .power_up = "low";

dffeas \epcs_slave_select_reg[14] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[14]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[14]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[14] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[14] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[14]~20 (
	.dataa(\p1_data_to_cpu[15]~14_combout ),
	.datab(\endofpacketvalue_reg[14]~q ),
	.datac(\epcs_slave_select_reg[14]~q ),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[14]~20_combout ),
	.cout());
defparam \p1_data_to_cpu[14]~20 .lut_mask = 16'hFAFC;
defparam \p1_data_to_cpu[14]~20 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[15] (
	.clk(clk),
	.d(data_from_cpu[15]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[15]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[15] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[15] .power_up = "low";

dffeas \epcs_slave_select_holding_reg[15] (
	.clk(clk),
	.d(data_from_cpu[15]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[15]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[15] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[15] .power_up = "low";

dffeas \epcs_slave_select_reg[15] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[15]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[15]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[15] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[15] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[15]~21 (
	.dataa(\p1_data_to_cpu[15]~14_combout ),
	.datab(\endofpacketvalue_reg[15]~q ),
	.datac(\epcs_slave_select_reg[15]~q ),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[15]~21_combout ),
	.cout());
defparam \p1_data_to_cpu[15]~21 .lut_mask = 16'hFAFC;
defparam \p1_data_to_cpu[15]~21 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[10] (
	.clk(clk),
	.d(data_from_cpu[10]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[10]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[10] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[10] .power_up = "low";

dffeas \epcs_slave_select_holding_reg[10] (
	.clk(clk),
	.d(data_from_cpu[10]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[10]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[10] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[10] .power_up = "low";

dffeas \epcs_slave_select_reg[10] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[10]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[10]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[10] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[10] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[10]~22 (
	.dataa(\endofpacketvalue_reg[10]~q ),
	.datab(\epcs_slave_select_reg[10]~q ),
	.datac(gnd),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[10]~22_combout ),
	.cout());
defparam \p1_data_to_cpu[10]~22 .lut_mask = 16'hAACC;
defparam \p1_data_to_cpu[10]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[10]~23 (
	.dataa(src_data_40),
	.datab(\p1_data_to_cpu[10]~22_combout ),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[10]~23_combout ),
	.cout());
defparam \p1_data_to_cpu[10]~23 .lut_mask = 16'hEFFE;
defparam \p1_data_to_cpu[10]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[10]~24 (
	.dataa(\p1_data_to_cpu[10]~23_combout ),
	.datab(\SSO_reg~q ),
	.datac(\p1_data_wr_strobe~0_combout ),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\p1_data_to_cpu[10]~24_combout ),
	.cout());
defparam \p1_data_to_cpu[10]~24 .lut_mask = 16'hFFFE;
defparam \p1_data_to_cpu[10]~24 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[9] (
	.clk(clk),
	.d(data_from_cpu[9]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[9]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[9] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[9] .power_up = "low";

dffeas \epcs_slave_select_holding_reg[9] (
	.clk(clk),
	.d(data_from_cpu[9]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[9]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[9] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[9] .power_up = "low";

dffeas \epcs_slave_select_reg[9] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[9]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[9]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[9] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[9] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[9]~25 (
	.dataa(src_data_38),
	.datab(\epcs_slave_select_reg[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p1_data_to_cpu[9]~25_combout ),
	.cout());
defparam \p1_data_to_cpu[9]~25 .lut_mask = 16'hEEEE;
defparam \p1_data_to_cpu[9]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_to_cpu[8]~3 (
	.dataa(src_data_40),
	.datab(gnd),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\data_to_cpu[8]~3_combout ),
	.cout());
defparam \data_to_cpu[8]~3 .lut_mask = 16'hAFFF;
defparam \data_to_cpu[8]~3 .sum_lutc_input = "datac";

dffeas iEOP_reg(
	.clk(clk),
	.d(data_from_cpu[9]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\iEOP_reg~q ),
	.prn(vcc));
defparam iEOP_reg.is_wysiwyg = "true";
defparam iEOP_reg.power_up = "low";

cycloneive_lcell_comb \EOP~0 (
	.dataa(\endofpacketvalue_reg[13]~q ),
	.datab(\endofpacketvalue_reg[12]~q ),
	.datac(\endofpacketvalue_reg[15]~q ),
	.datad(\endofpacketvalue_reg[14]~q ),
	.cin(gnd),
	.combout(\EOP~0_combout ),
	.cout());
defparam \EOP~0 .lut_mask = 16'h7FFF;
defparam \EOP~0 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[8] (
	.clk(clk),
	.d(data_from_cpu[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[8]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[8] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[8] .power_up = "low";

cycloneive_lcell_comb \EOP~1 (
	.dataa(\endofpacketvalue_reg[11]~q ),
	.datab(\endofpacketvalue_reg[9]~q ),
	.datac(\endofpacketvalue_reg[10]~q ),
	.datad(\endofpacketvalue_reg[8]~q ),
	.cin(gnd),
	.combout(\EOP~1_combout ),
	.cout());
defparam \EOP~1 .lut_mask = 16'h7FFF;
defparam \EOP~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~2 (
	.dataa(\rx_holding_reg[0]~q ),
	.datab(\rx_holding_reg[1]~q ),
	.datac(\endofpacketvalue_reg[1]~q ),
	.datad(\endofpacketvalue_reg[0]~q ),
	.cin(gnd),
	.combout(\EOP~2_combout ),
	.cout());
defparam \EOP~2 .lut_mask = 16'h6996;
defparam \EOP~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~3 (
	.dataa(\rx_holding_reg[2]~q ),
	.datab(\endofpacketvalue_reg[3]~q ),
	.datac(\rx_holding_reg[3]~q ),
	.datad(\endofpacketvalue_reg[2]~q ),
	.cin(gnd),
	.combout(\EOP~3_combout ),
	.cout());
defparam \EOP~3 .lut_mask = 16'h6996;
defparam \EOP~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~4 (
	.dataa(\endofpacketvalue_reg[4]~q ),
	.datab(\rx_holding_reg[5]~q ),
	.datac(\endofpacketvalue_reg[5]~q ),
	.datad(\rx_holding_reg[4]~q ),
	.cin(gnd),
	.combout(\EOP~4_combout ),
	.cout());
defparam \EOP~4 .lut_mask = 16'h6996;
defparam \EOP~4 .sum_lutc_input = "datac";

dffeas \endofpacketvalue_reg[7] (
	.clk(clk),
	.d(data_from_cpu[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[7]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[7] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[7] .power_up = "low";

dffeas \endofpacketvalue_reg[6] (
	.clk(clk),
	.d(data_from_cpu[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\endofpacketvalue_wr_strobe~combout ),
	.q(\endofpacketvalue_reg[6]~q ),
	.prn(vcc));
defparam \endofpacketvalue_reg[6] .is_wysiwyg = "true";
defparam \endofpacketvalue_reg[6] .power_up = "low";

dffeas \rx_holding_reg[6] (
	.clk(clk),
	.d(\shift_reg[6]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_holding_reg[3]~0_combout ),
	.q(\rx_holding_reg[6]~q ),
	.prn(vcc));
defparam \rx_holding_reg[6] .is_wysiwyg = "true";
defparam \rx_holding_reg[6] .power_up = "low";

dffeas \rx_holding_reg[7] (
	.clk(clk),
	.d(shift_reg_7),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_holding_reg[3]~0_combout ),
	.q(\rx_holding_reg[7]~q ),
	.prn(vcc));
defparam \rx_holding_reg[7] .is_wysiwyg = "true";
defparam \rx_holding_reg[7] .power_up = "low";

cycloneive_lcell_comb \EOP~5 (
	.dataa(\endofpacketvalue_reg[7]~q ),
	.datab(\endofpacketvalue_reg[6]~q ),
	.datac(\rx_holding_reg[6]~q ),
	.datad(\rx_holding_reg[7]~q ),
	.cin(gnd),
	.combout(\EOP~5_combout ),
	.cout());
defparam \EOP~5 .lut_mask = 16'h6996;
defparam \EOP~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~6 (
	.dataa(\EOP~2_combout ),
	.datab(\EOP~3_combout ),
	.datac(\EOP~4_combout ),
	.datad(\EOP~5_combout ),
	.cin(gnd),
	.combout(\EOP~6_combout ),
	.cout());
defparam \EOP~6 .lut_mask = 16'hFFFE;
defparam \EOP~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~7 (
	.dataa(data_from_cpu[7]),
	.datab(data_from_cpu[6]),
	.datac(\endofpacketvalue_reg[6]~q ),
	.datad(\endofpacketvalue_reg[7]~q ),
	.cin(gnd),
	.combout(\EOP~7_combout ),
	.cout());
defparam \EOP~7 .lut_mask = 16'h6996;
defparam \EOP~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~8 (
	.dataa(\EOP~0_combout ),
	.datab(\EOP~1_combout ),
	.datac(\EOP~6_combout ),
	.datad(\EOP~7_combout ),
	.cin(gnd),
	.combout(\EOP~8_combout ),
	.cout());
defparam \EOP~8 .lut_mask = 16'hFFFE;
defparam \EOP~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~9 (
	.dataa(data_from_cpu[5]),
	.datab(data_from_cpu[4]),
	.datac(\endofpacketvalue_reg[4]~q ),
	.datad(\endofpacketvalue_reg[5]~q ),
	.cin(gnd),
	.combout(\EOP~9_combout ),
	.cout());
defparam \EOP~9 .lut_mask = 16'h6996;
defparam \EOP~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~10 (
	.dataa(data_from_cpu[0]),
	.datab(data_from_cpu[1]),
	.datac(\endofpacketvalue_reg[1]~q ),
	.datad(\endofpacketvalue_reg[0]~q ),
	.cin(gnd),
	.combout(\EOP~10_combout ),
	.cout());
defparam \EOP~10 .lut_mask = 16'h6996;
defparam \EOP~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~11 (
	.dataa(data_from_cpu[3]),
	.datab(data_from_cpu[2]),
	.datac(\endofpacketvalue_reg[2]~q ),
	.datad(\endofpacketvalue_reg[3]~q ),
	.cin(gnd),
	.combout(\EOP~11_combout ),
	.cout());
defparam \EOP~11 .lut_mask = 16'h6996;
defparam \EOP~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~12 (
	.dataa(\EOP~10_combout ),
	.datab(\EOP~11_combout ),
	.datac(\EOP~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\EOP~12_combout ),
	.cout());
defparam \EOP~12 .lut_mask = 16'hFEFE;
defparam \EOP~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~13 (
	.dataa(\p1_rd_strobe~0_combout ),
	.datab(\p1_data_rd_strobe~0_combout ),
	.datac(\EOP~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\EOP~13_combout ),
	.cout());
defparam \EOP~13 .lut_mask = 16'hFEFE;
defparam \EOP~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~14 (
	.dataa(\EOP~9_combout ),
	.datab(\p1_data_wr_strobe~combout ),
	.datac(\EOP~12_combout ),
	.datad(\EOP~13_combout ),
	.cin(gnd),
	.combout(\EOP~14_combout ),
	.cout());
defparam \EOP~14 .lut_mask = 16'hFFFE;
defparam \EOP~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \EOP~15 (
	.dataa(\EOP~q ),
	.datab(\status_wr_strobe~combout ),
	.datac(\EOP~8_combout ),
	.datad(\EOP~14_combout ),
	.cin(gnd),
	.combout(\EOP~15_combout ),
	.cout());
defparam \EOP~15 .lut_mask = 16'hFFFB;
defparam \EOP~15 .sum_lutc_input = "datac";

dffeas EOP(
	.clk(clk),
	.d(\EOP~15_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\EOP~q ),
	.prn(vcc));
defparam EOP.is_wysiwyg = "true";
defparam EOP.power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[9]~26 (
	.dataa(\iEOP_reg~q ),
	.datab(\EOP~q ),
	.datac(src_data_40),
	.datad(\data_to_cpu[4]~2_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[9]~26_combout ),
	.cout());
defparam \p1_data_to_cpu[9]~26 .lut_mask = 16'hEFFE;
defparam \p1_data_to_cpu[9]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[9]~27 (
	.dataa(\endofpacketvalue_reg[9]~q ),
	.datab(\p1_data_to_cpu[9]~25_combout ),
	.datac(\data_to_cpu[8]~3_combout ),
	.datad(\p1_data_to_cpu[9]~26_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[9]~27_combout ),
	.cout());
defparam \p1_data_to_cpu[9]~27 .lut_mask = 16'hEFFE;
defparam \p1_data_to_cpu[9]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[9]~28 (
	.dataa(\p1_data_to_cpu[9]~27_combout ),
	.datab(src_data_40),
	.datac(src_data_39),
	.datad(gnd),
	.cin(gnd),
	.combout(\p1_data_to_cpu[9]~28_combout ),
	.cout());
defparam \p1_data_to_cpu[9]~28 .lut_mask = 16'hFEFE;
defparam \p1_data_to_cpu[9]~28 .sum_lutc_input = "datac";

dffeas \epcs_slave_select_holding_reg[8] (
	.clk(clk),
	.d(data_from_cpu[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[8]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[8] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[8] .power_up = "low";

dffeas \epcs_slave_select_reg[8] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[8]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[8]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[8] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[8] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[8]~29 (
	.dataa(src_data_38),
	.datab(\epcs_slave_select_reg[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p1_data_to_cpu[8]~29_combout ),
	.cout());
defparam \p1_data_to_cpu[8]~29 .lut_mask = 16'hEEEE;
defparam \p1_data_to_cpu[8]~29 .sum_lutc_input = "datac";

dffeas iE_reg(
	.clk(clk),
	.d(data_from_cpu[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\iE_reg~q ),
	.prn(vcc));
defparam iE_reg.is_wysiwyg = "true";
defparam iE_reg.power_up = "low";

cycloneive_lcell_comb E(
	.dataa(\TOE~q ),
	.datab(\ROE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E~combout ),
	.cout());
defparam E.lut_mask = 16'hEEEE;
defparam E.sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[8]~30 (
	.dataa(\iE_reg~q ),
	.datab(\E~combout ),
	.datac(src_data_40),
	.datad(\data_to_cpu[4]~2_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[8]~30_combout ),
	.cout());
defparam \p1_data_to_cpu[8]~30 .lut_mask = 16'hEFFE;
defparam \p1_data_to_cpu[8]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[8]~31 (
	.dataa(\endofpacketvalue_reg[8]~q ),
	.datab(\p1_data_to_cpu[8]~29_combout ),
	.datac(\data_to_cpu[8]~3_combout ),
	.datad(\p1_data_to_cpu[8]~30_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[8]~31_combout ),
	.cout());
defparam \p1_data_to_cpu[8]~31 .lut_mask = 16'hEFFE;
defparam \p1_data_to_cpu[8]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[8]~32 (
	.dataa(\p1_data_to_cpu[8]~31_combout ),
	.datab(src_data_40),
	.datac(src_data_39),
	.datad(gnd),
	.cin(gnd),
	.combout(\p1_data_to_cpu[8]~32_combout ),
	.cout());
defparam \p1_data_to_cpu[8]~32 .lut_mask = 16'hFEFE;
defparam \p1_data_to_cpu[8]~32 .sum_lutc_input = "datac";

dffeas iRRDY_reg(
	.clk(clk),
	.d(data_from_cpu[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\iRRDY_reg~q ),
	.prn(vcc));
defparam iRRDY_reg.is_wysiwyg = "true";
defparam iRRDY_reg.power_up = "low";

dffeas \epcs_slave_select_holding_reg[7] (
	.clk(clk),
	.d(data_from_cpu[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[7]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[7] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[7] .power_up = "low";

dffeas \epcs_slave_select_reg[7] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[7]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[7]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[7] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[7] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[7]~33 (
	.dataa(\data_to_cpu[4]~2_combout ),
	.datab(\epcs_slave_select_reg[7]~q ),
	.datac(src_data_40),
	.datad(\RRDY~q ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[7]~33_combout ),
	.cout());
defparam \p1_data_to_cpu[7]~33 .lut_mask = 16'hFFDE;
defparam \p1_data_to_cpu[7]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[7]~34 (
	.dataa(\iRRDY_reg~q ),
	.datab(\data_to_cpu[4]~2_combout ),
	.datac(\p1_data_to_cpu[7]~33_combout ),
	.datad(\endofpacketvalue_reg[7]~q ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[7]~34_combout ),
	.cout());
defparam \p1_data_to_cpu[7]~34 .lut_mask = 16'hFFBE;
defparam \p1_data_to_cpu[7]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[7]~35 (
	.dataa(\p1_data_to_cpu[7]~34_combout ),
	.datab(\rx_holding_reg[7]~q ),
	.datac(gnd),
	.datad(\data_to_cpu[0]~1_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[7]~35_combout ),
	.cout());
defparam \p1_data_to_cpu[7]~35 .lut_mask = 16'hAACC;
defparam \p1_data_to_cpu[7]~35 .sum_lutc_input = "datac";

dffeas iTRDY_reg(
	.clk(clk),
	.d(data_from_cpu[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\iTRDY_reg~q ),
	.prn(vcc));
defparam iTRDY_reg.is_wysiwyg = "true";
defparam iTRDY_reg.power_up = "low";

dffeas \epcs_slave_select_holding_reg[6] (
	.clk(clk),
	.d(data_from_cpu[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slaveselect_wr_strobe~0_combout ),
	.q(\epcs_slave_select_holding_reg[6]~q ),
	.prn(vcc));
defparam \epcs_slave_select_holding_reg[6] .is_wysiwyg = "true";
defparam \epcs_slave_select_holding_reg[6] .power_up = "low";

dffeas \epcs_slave_select_reg[6] (
	.clk(clk),
	.d(\epcs_slave_select_holding_reg[6]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\epcs_slave_select_reg[6]~q ),
	.prn(vcc));
defparam \epcs_slave_select_reg[6] .is_wysiwyg = "true";
defparam \epcs_slave_select_reg[6] .power_up = "low";

cycloneive_lcell_comb \p1_data_to_cpu[6]~36 (
	.dataa(\data_to_cpu[4]~2_combout ),
	.datab(\epcs_slave_select_reg[6]~q ),
	.datac(src_data_40),
	.datad(\TRDY~0_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[6]~36_combout ),
	.cout());
defparam \p1_data_to_cpu[6]~36 .lut_mask = 16'hDEFF;
defparam \p1_data_to_cpu[6]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[6]~37 (
	.dataa(\iTRDY_reg~q ),
	.datab(\data_to_cpu[4]~2_combout ),
	.datac(\p1_data_to_cpu[6]~36_combout ),
	.datad(\endofpacketvalue_reg[6]~q ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[6]~37_combout ),
	.cout());
defparam \p1_data_to_cpu[6]~37 .lut_mask = 16'hFFBE;
defparam \p1_data_to_cpu[6]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_data_to_cpu[6]~38 (
	.dataa(\p1_data_to_cpu[6]~37_combout ),
	.datab(\rx_holding_reg[6]~q ),
	.datac(gnd),
	.datad(\data_to_cpu[0]~1_combout ),
	.cin(gnd),
	.combout(\p1_data_to_cpu[6]~38_combout ),
	.cout());
defparam \p1_data_to_cpu[6]~38 .lut_mask = 16'hAACC;
defparam \p1_data_to_cpu[6]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \irq_reg~0 (
	.dataa(\iE_reg~q ),
	.datab(\TOE~q ),
	.datac(\iTOE_reg~q ),
	.datad(\ROE~q ),
	.cin(gnd),
	.combout(\irq_reg~0_combout ),
	.cout());
defparam \irq_reg~0 .lut_mask = 16'hFFFE;
defparam \irq_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \irq_reg~1 (
	.dataa(\iEOP_reg~q ),
	.datab(\iRRDY_reg~q ),
	.datac(\RRDY~q ),
	.datad(\EOP~q ),
	.cin(gnd),
	.combout(\irq_reg~1_combout ),
	.cout());
defparam \irq_reg~1 .lut_mask = 16'hFFFE;
defparam \irq_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \irq_reg~2 (
	.dataa(\iROE_reg~q ),
	.datab(\ROE~q ),
	.datac(\iTRDY_reg~q ),
	.datad(\TRDY~0_combout ),
	.cin(gnd),
	.combout(\irq_reg~2_combout ),
	.cout());
defparam \irq_reg~2 .lut_mask = 16'hFEFF;
defparam \irq_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \irq_reg~3 (
	.dataa(\irq_reg~0_combout ),
	.datab(\irq_reg~1_combout ),
	.datac(\irq_reg~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\irq_reg~3_combout ),
	.cout());
defparam \irq_reg~3 .lut_mask = 16'hFEFE;
defparam \irq_reg~3 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_jtag (
	tdo,
	altera_reset_synchronizer_int_chain_out,
	rst1,
	b_full,
	out_data_toggle_flopped,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	dreg_0,
	av_waitrequest1,
	mem_used_1,
	out_data_buffer_66,
	out_data_buffer_38,
	out_data_buffer_7,
	out_data_buffer_65,
	out_data_buffer_0,
	b_full1,
	counter_reg_bit_21,
	counter_reg_bit_11,
	counter_reg_bit_51,
	counter_reg_bit_41,
	counter_reg_bit_31,
	counter_reg_bit_01,
	out_data_buffer_1,
	read_01,
	av_readdata_0,
	av_readdata_9,
	av_irq1,
	av_readdata_1,
	av_readdata_2,
	av_readdata_3,
	av_readdata_4,
	av_readdata_5,
	av_readdata_6,
	av_readdata_7,
	out_data_buffer_2,
	rvalid1,
	woverflow1,
	ac1,
	av_readdata_8,
	out_data_buffer_3,
	out_data_buffer_10,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	tdo;
input 	altera_reset_synchronizer_int_chain_out;
output 	rst1;
output 	b_full;
input 	out_data_toggle_flopped;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	dreg_0;
output 	av_waitrequest1;
input 	mem_used_1;
input 	out_data_buffer_66;
input 	out_data_buffer_38;
input 	out_data_buffer_7;
input 	out_data_buffer_65;
input 	out_data_buffer_0;
output 	b_full1;
output 	counter_reg_bit_21;
output 	counter_reg_bit_11;
output 	counter_reg_bit_51;
output 	counter_reg_bit_41;
output 	counter_reg_bit_31;
output 	counter_reg_bit_01;
input 	out_data_buffer_1;
output 	read_01;
output 	av_readdata_0;
output 	av_readdata_9;
output 	av_irq1;
output 	av_readdata_1;
output 	av_readdata_2;
output 	av_readdata_3;
output 	av_readdata_4;
output 	av_readdata_5;
output 	av_readdata_6;
output 	av_readdata_7;
input 	out_data_buffer_2;
output 	rvalid1;
output 	woverflow1;
output 	ac1;
output 	av_readdata_8;
input 	out_data_buffer_3;
input 	out_data_buffer_10;
input 	out_data_buffer_4;
input 	out_data_buffer_5;
input 	out_data_buffer_6;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \t_dav~q ;
wire \niosII_jtag_alt_jtag_atlantic|rvalid0~q ;
wire \r_val~q ;
wire \niosII_jtag_alt_jtag_atlantic|r_ena1~q ;
wire \niosII_jtag_alt_jtag_atlantic|t_ena~q ;
wire \the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \fifo_wr~q ;
wire \wr_rfifo~combout ;
wire \fifo_wr~0_combout ;
wire \niosII_jtag_alt_jtag_atlantic|wdata[0]~q ;
wire \niosII_jtag_alt_jtag_atlantic|t_pause~q ;
wire \niosII_jtag_alt_jtag_atlantic|wdata[1]~q ;
wire \niosII_jtag_alt_jtag_atlantic|wdata[2]~q ;
wire \niosII_jtag_alt_jtag_atlantic|wdata[3]~q ;
wire \niosII_jtag_alt_jtag_atlantic|wdata[4]~q ;
wire \niosII_jtag_alt_jtag_atlantic|wdata[5]~q ;
wire \niosII_jtag_alt_jtag_atlantic|wdata[6]~q ;
wire \niosII_jtag_alt_jtag_atlantic|wdata[7]~q ;
wire \fifo_rd~0_combout ;
wire \av_waitrequest~0_combout ;
wire \fifo_rd~2_combout ;
wire \ien_AF~0_combout ;
wire \ien_AF~q ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \ien_AE~q ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \Add0~0_combout ;
wire \Add0~2_combout ;
wire \LessThan1~0_combout ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \LessThan1~1_combout ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \LessThan1~2_combout ;
wire \fifo_AF~q ;
wire \fifo_rd~1_combout ;
wire \rvalid~0_combout ;
wire \fifo_wr~1_combout ;
wire \woverflow~0_combout ;
wire \ac~0_combout ;
wire \ac~1_combout ;


niosII_niosII_jtag_scfifo_w the_niosII_jtag_scfifo_w(
	.q_b_7(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_0(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_non_empty(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val(\r_val~0_combout ),
	.fifo_wr(\fifo_wr~q ),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_0(out_data_buffer_0),
	.b_full(b_full1),
	.counter_reg_bit_2(counter_reg_bit_21),
	.counter_reg_bit_1(counter_reg_bit_11),
	.counter_reg_bit_5(counter_reg_bit_51),
	.counter_reg_bit_4(counter_reg_bit_41),
	.counter_reg_bit_3(counter_reg_bit_31),
	.counter_reg_bit_0(counter_reg_bit_01),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_6(out_data_buffer_6),
	.clk_clk(clk_clk));

niosII_niosII_jtag_scfifo_r the_niosII_jtag_scfifo_r(
	.q_b_0(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(\niosII_jtag_alt_jtag_atlantic|t_ena~q ),
	.fifo_rd(\fifo_rd~1_combout ),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_0(\niosII_jtag_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\niosII_jtag_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\niosII_jtag_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\niosII_jtag_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\niosII_jtag_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\niosII_jtag_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\niosII_jtag_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\niosII_jtag_alt_jtag_atlantic|wdata[7]~q ),
	.clk_clk(clk_clk));

niosII_alt_jtag_atlantic niosII_jtag_alt_jtag_atlantic(
	.r_dat({\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ,\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ,\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ,
\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ,\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ,\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ,
\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ,\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.tdo1(tdo),
	.rst_n(altera_reset_synchronizer_int_chain_out),
	.rst11(rst1),
	.t_dav(\t_dav~q ),
	.rvalid01(\niosII_jtag_alt_jtag_atlantic|rvalid0~q ),
	.r_val(\r_val~q ),
	.r_ena11(\niosII_jtag_alt_jtag_atlantic|r_ena1~q ),
	.t_ena1(\niosII_jtag_alt_jtag_atlantic|t_ena~q ),
	.wdata_0(\niosII_jtag_alt_jtag_atlantic|wdata[0]~q ),
	.t_pause1(\niosII_jtag_alt_jtag_atlantic|t_pause~q ),
	.wdata_1(\niosII_jtag_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\niosII_jtag_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\niosII_jtag_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\niosII_jtag_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\niosII_jtag_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\niosII_jtag_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\niosII_jtag_alt_jtag_atlantic|wdata[7]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

cycloneive_lcell_comb \r_val~0 (
	.dataa(\the_niosII_jtag_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datab(\r_val~q ),
	.datac(\niosII_jtag_alt_jtag_atlantic|r_ena1~q ),
	.datad(\niosII_jtag_alt_jtag_atlantic|rvalid0~q ),
	.cin(gnd),
	.combout(\r_val~0_combout ),
	.cout());
defparam \r_val~0 .lut_mask = 16'hBFFF;
defparam \r_val~0 .sum_lutc_input = "datac";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cycloneive_lcell_comb wr_rfifo(
	.dataa(\niosII_jtag_alt_jtag_atlantic|t_ena~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(b_full),
	.cin(gnd),
	.combout(\wr_rfifo~combout ),
	.cout());
defparam wr_rfifo.lut_mask = 16'hAAFF;
defparam wr_rfifo.sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_wr~0 (
	.dataa(out_data_buffer_38),
	.datab(b_full1),
	.datac(\fifo_rd~0_combout ),
	.datad(out_data_buffer_65),
	.cin(gnd),
	.combout(\fifo_wr~0_combout ),
	.cout());
defparam \fifo_wr~0 .lut_mask = 16'hFFF7;
defparam \fifo_wr~0 .sum_lutc_input = "datac";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\av_waitrequest~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest1),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

cycloneive_lcell_comb \av_readdata[0]~0 (
	.dataa(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\ien_AF~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_0),
	.cout());
defparam \av_readdata[0]~0 .lut_mask = 16'hAACC;
defparam \av_readdata[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[9] (
	.dataa(\fifo_AE~q ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_9),
	.cout());
defparam \av_readdata[9] .lut_mask = 16'hEEEE;
defparam \av_readdata[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb av_irq(
	.dataa(av_readdata_9),
	.datab(\ien_AF~q ),
	.datac(\pause_irq~q ),
	.datad(\fifo_AF~q ),
	.cin(gnd),
	.combout(av_irq1),
	.cout());
defparam av_irq.lut_mask = 16'hFFFE;
defparam av_irq.sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[1]~1 (
	.dataa(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_1),
	.cout());
defparam \av_readdata[1]~1 .lut_mask = 16'hAACC;
defparam \av_readdata[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[2]~2 (
	.dataa(read_01),
	.datab(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_2),
	.cout());
defparam \av_readdata[2]~2 .lut_mask = 16'hEEEE;
defparam \av_readdata[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[3]~3 (
	.dataa(read_01),
	.datab(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_3),
	.cout());
defparam \av_readdata[3]~3 .lut_mask = 16'hEEEE;
defparam \av_readdata[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[4]~4 (
	.dataa(read_01),
	.datab(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_4),
	.cout());
defparam \av_readdata[4]~4 .lut_mask = 16'hEEEE;
defparam \av_readdata[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[5]~5 (
	.dataa(read_01),
	.datab(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_5),
	.cout());
defparam \av_readdata[5]~5 .lut_mask = 16'hEEEE;
defparam \av_readdata[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[6]~6 (
	.dataa(read_01),
	.datab(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_6),
	.cout());
defparam \av_readdata[6]~6 .lut_mask = 16'hEEEE;
defparam \av_readdata[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[7]~7 (
	.dataa(read_01),
	.datab(\the_niosII_jtag_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_7),
	.cout());
defparam \av_readdata[7]~7 .lut_mask = 16'hEEEE;
defparam \av_readdata[7]~7 .sum_lutc_input = "datac";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

cycloneive_lcell_comb \av_readdata[8]~8 (
	.dataa(\ien_AF~q ),
	.datab(\pause_irq~q ),
	.datac(\fifo_AF~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_8),
	.cout());
defparam \av_readdata[8]~8 .lut_mask = 16'hFEFE;
defparam \av_readdata[8]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_rd~0 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(av_waitrequest1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\fifo_rd~0_combout ),
	.cout());
defparam \fifo_rd~0 .lut_mask = 16'h6FFF;
defparam \fifo_rd~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest~0 (
	.dataa(\fifo_rd~0_combout ),
	.datab(out_data_buffer_66),
	.datac(out_data_buffer_65),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_waitrequest~0_combout ),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hFEFE;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_rd~2 (
	.dataa(\fifo_rd~0_combout ),
	.datab(out_data_buffer_66),
	.datac(gnd),
	.datad(out_data_buffer_38),
	.cin(gnd),
	.combout(\fifo_rd~2_combout ),
	.cout());
defparam \fifo_rd~2 .lut_mask = 16'hEEFF;
defparam \fifo_rd~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ien_AF~0 (
	.dataa(\fifo_rd~0_combout ),
	.datab(out_data_buffer_38),
	.datac(out_data_buffer_65),
	.datad(gnd),
	.cin(gnd),
	.combout(\ien_AF~0_combout ),
	.cout());
defparam \ien_AF~0 .lut_mask = 16'hFEFE;
defparam \ien_AF~0 .sum_lutc_input = "datac";

dffeas ien_AF(
	.clk(clk_clk),
	.d(out_data_buffer_0),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AF~0_combout ),
	.q(\ien_AF~q ),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

cycloneive_lcell_comb \LessThan0~0 (
	.dataa(counter_reg_bit_31),
	.datab(counter_reg_bit_21),
	.datac(counter_reg_bit_11),
	.datad(counter_reg_bit_01),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'hFFFE;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~1 (
	.dataa(b_full1),
	.datab(counter_reg_bit_51),
	.datac(counter_reg_bit_41),
	.datad(\LessThan0~0_combout ),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

dffeas ien_AE(
	.clk(clk_clk),
	.d(out_data_buffer_1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AF~0_combout ),
	.q(\ien_AE~q ),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

cycloneive_lcell_comb \pause_irq~0 (
	.dataa(b_non_empty),
	.datab(\niosII_jtag_alt_jtag_atlantic|t_pause~q ),
	.datac(\pause_irq~q ),
	.datad(read_01),
	.cin(gnd),
	.combout(\pause_irq~0_combout ),
	.cout());
defparam \pause_irq~0 .lut_mask = 16'hFEFF;
defparam \pause_irq~0 .sum_lutc_input = "datac";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(counter_reg_bit_0),
	.datab(counter_reg_bit_1),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h6677;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~2 (
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5AAF;
defparam \Add0~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~4 (
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5A5F;
defparam \Add0~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~0 (
	.dataa(\Add0~4_combout ),
	.datab(counter_reg_bit_0),
	.datac(\Add0~0_combout ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\LessThan1~0_combout ),
	.cout());
defparam \LessThan1~0 .lut_mask = 16'hFFFE;
defparam \LessThan1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~6 (
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5AAF;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~8 (
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5A5F;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~1 (
	.dataa(\Add0~6_combout ),
	.datab(\Add0~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan1~1_combout ),
	.cout());
defparam \LessThan1~1 .lut_mask = 16'hEEEE;
defparam \LessThan1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~10 (
	.dataa(b_full),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5AAF;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout());
defparam \Add0~12 .lut_mask = 16'hF0F0;
defparam \Add0~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~2 (
	.dataa(\LessThan1~0_combout ),
	.datab(\LessThan1~1_combout ),
	.datac(\Add0~10_combout ),
	.datad(\Add0~12_combout ),
	.cin(gnd),
	.combout(\LessThan1~2_combout ),
	.cout());
defparam \LessThan1~2 .lut_mask = 16'h7FFF;
defparam \LessThan1~2 .sum_lutc_input = "datac";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cycloneive_lcell_comb \fifo_rd~1 (
	.dataa(b_non_empty),
	.datab(\fifo_rd~0_combout ),
	.datac(out_data_buffer_66),
	.datad(out_data_buffer_38),
	.cin(gnd),
	.combout(\fifo_rd~1_combout ),
	.cout());
defparam \fifo_rd~1 .lut_mask = 16'hFEFF;
defparam \fifo_rd~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rvalid~0 (
	.dataa(\fifo_rd~1_combout ),
	.datab(rvalid1),
	.datac(gnd),
	.datad(\fifo_rd~2_combout ),
	.cin(gnd),
	.combout(\rvalid~0_combout ),
	.cout());
defparam \rvalid~0 .lut_mask = 16'hEEFF;
defparam \rvalid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_wr~1 (
	.dataa(\fifo_rd~0_combout ),
	.datab(out_data_buffer_65),
	.datac(gnd),
	.datad(out_data_buffer_38),
	.cin(gnd),
	.combout(\fifo_wr~1_combout ),
	.cout());
defparam \fifo_wr~1 .lut_mask = 16'hEEFF;
defparam \fifo_wr~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \woverflow~0 (
	.dataa(b_full1),
	.datab(woverflow1),
	.datac(gnd),
	.datad(\fifo_wr~1_combout ),
	.cin(gnd),
	.combout(\woverflow~0_combout ),
	.cout());
defparam \woverflow~0 .lut_mask = 16'hAACC;
defparam \woverflow~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ac~0 (
	.dataa(\niosII_jtag_alt_jtag_atlantic|t_ena~q ),
	.datab(\niosII_jtag_alt_jtag_atlantic|t_pause~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac~0_combout ),
	.cout());
defparam \ac~0 .lut_mask = 16'hEEEE;
defparam \ac~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ac~1 (
	.dataa(\ac~0_combout ),
	.datab(ac1),
	.datac(\ien_AF~0_combout ),
	.datad(out_data_buffer_10),
	.cin(gnd),
	.combout(\ac~1_combout ),
	.cout());
defparam \ac~1 .lut_mask = 16'hEFFF;
defparam \ac~1 .sum_lutc_input = "datac";

endmodule

module niosII_alt_jtag_atlantic (
	r_dat,
	tdo1,
	rst_n,
	rst11,
	t_dav,
	rvalid01,
	r_val,
	r_ena11,
	t_ena1,
	wdata_0,
	t_pause1,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	tdo1;
input 	rst_n;
output 	rst11;
input 	t_dav;
output 	rvalid01;
input 	r_val;
output 	r_ena11;
output 	t_ena1;
output 	wdata_0;
output 	t_pause1;
output 	wdata_1;
output 	wdata_2;
output 	wdata_3;
output 	wdata_4;
output 	wdata_5;
output 	wdata_6;
output 	wdata_7;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \state~1_combout ;
wire \always0~0_combout ;
wire \state~0_combout ;
wire \state~2_combout ;
wire \state~q ;
wire \count~9_combout ;
wire \td_shift[0]~4_combout ;
wire \count[2]~q ;
wire \count~8_combout ;
wire \count[3]~q ;
wire \count~7_combout ;
wire \count[4]~q ;
wire \count~6_combout ;
wire \count[5]~q ;
wire \count~5_combout ;
wire \count[6]~q ;
wire \count~4_combout ;
wire \count[7]~q ;
wire \count~2_combout ;
wire \count[8]~q ;
wire \count[9]~0_combout ;
wire \count[9]~q ;
wire \count~3_combout ;
wire \count[0]~q ;
wire \count~1_combout ;
wire \count[1]~q ;
wire \write~2_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift~10_combout ;
wire \td_shift[10]~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~7_combout ;
wire \td_shift[9]~q ;
wire \td_shift~1_combout ;
wire \rdata[6]~q ;
wire \td_shift~21_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~19_combout ;
wire \td_shift~20_combout ;
wire \td_shift[7]~q ;
wire \rdata[4]~q ;
wire \td_shift~17_combout ;
wire \td_shift~18_combout ;
wire \td_shift[6]~q ;
wire \rdata[3]~q ;
wire \td_shift~15_combout ;
wire \td_shift~16_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~13_combout ;
wire \td_shift~14_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~11_combout ;
wire \td_shift~12_combout ;
wire \td_shift[3]~q ;
wire \rdata[0]~q ;
wire \td_shift~8_combout ;
wire \td_shift~9_combout ;
wire \td_shift[2]~q ;
wire \write_stalled~2_combout ;
wire \write_stalled~4_combout ;
wire \write_stalled~3_combout ;
wire \write_stalled~q ;
wire \td_shift~5_combout ;
wire \td_shift~6_combout ;
wire \td_shift[1]~q ;
wire \rvalid~q ;
wire \td_shift~0_combout ;
wire \td_shift~2_combout ;
wire \td_shift~3_combout ;
wire \td_shift[0]~q ;
wire \rvalid0~0_combout ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \read_req~q ;
wire \rvalid0~1_combout ;
wire \rst2~q ;
wire \rvalid0~2_combout ;
wire \write~4_combout ;
wire \write~3_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \write_valid~q ;
wire \t_ena~2_combout ;
wire \t_ena~3_combout ;
wire \always2~0_combout ;
wire \t_pause~0_combout ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \t_pause~1_combout ;


dffeas tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tdo1),
	.prn(vcc));
defparam tdo.is_wysiwyg = "true";
defparam tdo.power_up = "low";

dffeas rst1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rst11),
	.prn(vcc));
defparam rst1.is_wysiwyg = "true";
defparam rst1.power_up = "low";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid01),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_ena11),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

dffeas t_ena(
	.clk(clk),
	.d(\t_ena~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena1),
	.prn(vcc));
defparam t_ena.is_wysiwyg = "true";
defparam t_ena.power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas t_pause(
	.clk(clk),
	.d(\t_pause~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause1),
	.prn(vcc));
defparam t_pause.is_wysiwyg = "true";
defparam t_pause.power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~3_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~3_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~3_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~3_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~3_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~3_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~3_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

cycloneive_lcell_comb \tck_t_dav~0 (
	.dataa(t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tck_t_dav~0_combout ),
	.cout());
defparam \tck_t_dav~0 .lut_mask = 16'h5555;
defparam \tck_t_dav~0 .sum_lutc_input = "datac";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cycloneive_lcell_comb \state~1 (
	.dataa(\state~q ),
	.datab(virtual_ir_scan_reg),
	.datac(splitter_nodes_receive_0_3),
	.datad(state_3),
	.cin(gnd),
	.combout(\state~1_combout ),
	.cout());
defparam \state~1 .lut_mask = 16'hEFFF;
defparam \state~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(gnd),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hAAFF;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~0 (
	.dataa(altera_internal_jtag1),
	.datab(gnd),
	.datac(irf_reg_0_1),
	.datad(\state~q ),
	.cin(gnd),
	.combout(\state~0_combout ),
	.cout());
defparam \state~0 .lut_mask = 16'hAFFF;
defparam \state~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~2 (
	.dataa(\state~1_combout ),
	.datab(state_4),
	.datac(\always0~0_combout ),
	.datad(\state~0_combout ),
	.cin(gnd),
	.combout(\state~2_combout ),
	.cout());
defparam \state~2 .lut_mask = 16'hFFFE;
defparam \state~2 .sum_lutc_input = "datac";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cycloneive_lcell_comb \count~9 (
	.dataa(\count[1]~q ),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~9_combout ),
	.cout());
defparam \count~9 .lut_mask = 16'hEEEE;
defparam \count~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift[0]~4 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(state_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\td_shift[0]~4_combout ),
	.cout());
defparam \td_shift[0]~4 .lut_mask = 16'hFEFF;
defparam \td_shift[0]~4 .sum_lutc_input = "datac";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cycloneive_lcell_comb \count~8 (
	.dataa(state_4),
	.datab(\count[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~8_combout ),
	.cout());
defparam \count~8 .lut_mask = 16'hEEEE;
defparam \count~8 .sum_lutc_input = "datac";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cycloneive_lcell_comb \count~7 (
	.dataa(state_4),
	.datab(\count[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~7_combout ),
	.cout());
defparam \count~7 .lut_mask = 16'hEEEE;
defparam \count~7 .sum_lutc_input = "datac";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneive_lcell_comb \count~6 (
	.dataa(state_4),
	.datab(\count[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~6_combout ),
	.cout());
defparam \count~6 .lut_mask = 16'hEEEE;
defparam \count~6 .sum_lutc_input = "datac";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cycloneive_lcell_comb \count~5 (
	.dataa(state_4),
	.datab(\count[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~5_combout ),
	.cout());
defparam \count~5 .lut_mask = 16'hEEEE;
defparam \count~5 .sum_lutc_input = "datac";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneive_lcell_comb \count~4 (
	.dataa(state_4),
	.datab(\count[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~4_combout ),
	.cout());
defparam \count~4 .lut_mask = 16'hEEEE;
defparam \count~4 .sum_lutc_input = "datac";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count~4_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneive_lcell_comb \count~2 (
	.dataa(state_4),
	.datab(\count[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~2_combout ),
	.cout());
defparam \count~2 .lut_mask = 16'hEEEE;
defparam \count~2 .sum_lutc_input = "datac";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cycloneive_lcell_comb \count[9]~0 (
	.dataa(state_4),
	.datab(\state~0_combout ),
	.datac(\count[8]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[9]~0_combout ),
	.cout());
defparam \count[9]~0 .lut_mask = 16'h7F7F;
defparam \count[9]~0 .sum_lutc_input = "datac";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cycloneive_lcell_comb \count~3 (
	.dataa(state_4),
	.datab(gnd),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
defparam \count~3 .lut_mask = 16'hAAFF;
defparam \count~3 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneive_lcell_comb \count~1 (
	.dataa(state_4),
	.datab(\count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~1_combout ),
	.cout());
defparam \count~1 .lut_mask = 16'hEEEE;
defparam \count~1 .sum_lutc_input = "datac";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneive_lcell_comb \write~2 (
	.dataa(\state~q ),
	.datab(state_4),
	.datac(\always0~0_combout ),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\write~2_combout ),
	.cout());
defparam \write~2 .lut_mask = 16'hFEFF;
defparam \write~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \user_saw_rvalid~0 (
	.dataa(\td_shift[0]~q ),
	.datab(\user_saw_rvalid~q ),
	.datac(\count[0]~q ),
	.datad(\write~2_combout ),
	.cin(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.cout());
defparam \user_saw_rvalid~0 .lut_mask = 16'hEFFE;
defparam \user_saw_rvalid~0 .sum_lutc_input = "datac";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

cycloneive_lcell_comb \td_shift~10 (
	.dataa(altera_internal_jtag1),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~10_combout ),
	.cout());
defparam \td_shift~10 .lut_mask = 16'hEEEE;
defparam \td_shift~10 .sum_lutc_input = "datac";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

cycloneive_lcell_comb \r_ena~0 (
	.dataa(r_val),
	.datab(r_ena11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\r_ena~0_combout ),
	.cout());
defparam \r_ena~0 .lut_mask = 16'hEEEE;
defparam \r_ena~0 .sum_lutc_input = "datac";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cycloneive_lcell_comb \td_shift~7 (
	.dataa(\td_shift[10]~q ),
	.datab(\rdata[7]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~7_combout ),
	.cout());
defparam \td_shift~7 .lut_mask = 16'hAACC;
defparam \td_shift~7 .sum_lutc_input = "datac";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cycloneive_lcell_comb \td_shift~1 (
	.dataa(\state~q ),
	.datab(\count[1]~q ),
	.datac(\user_saw_rvalid~q ),
	.datad(\td_shift[9]~q ),
	.cin(gnd),
	.combout(\td_shift~1_combout ),
	.cout());
defparam \td_shift~1 .lut_mask = 16'hEFFF;
defparam \td_shift~1 .sum_lutc_input = "datac";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cycloneive_lcell_comb \td_shift~21 (
	.dataa(\td_shift[9]~q ),
	.datab(\rdata[6]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~21_combout ),
	.cout());
defparam \td_shift~21 .lut_mask = 16'hAACC;
defparam \td_shift~21 .sum_lutc_input = "datac";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~21_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cycloneive_lcell_comb \td_shift~19 (
	.dataa(\td_shift[8]~q ),
	.datab(\rdata[5]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~19_combout ),
	.cout());
defparam \td_shift~19 .lut_mask = 16'hACAC;
defparam \td_shift~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~20 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~1_combout ),
	.datad(\td_shift~19_combout ),
	.cin(gnd),
	.combout(\td_shift~20_combout ),
	.cout());
defparam \td_shift~20 .lut_mask = 16'hFFEF;
defparam \td_shift~20 .sum_lutc_input = "datac";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~20_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

cycloneive_lcell_comb \td_shift~17 (
	.dataa(\td_shift[7]~q ),
	.datab(\rdata[4]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~17_combout ),
	.cout());
defparam \td_shift~17 .lut_mask = 16'hAACC;
defparam \td_shift~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~18 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~17_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~18_combout ),
	.cout());
defparam \td_shift~18 .lut_mask = 16'hACFF;
defparam \td_shift~18 .sum_lutc_input = "datac";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~18_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

cycloneive_lcell_comb \td_shift~15 (
	.dataa(\td_shift[6]~q ),
	.datab(\rdata[3]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~15_combout ),
	.cout());
defparam \td_shift~15 .lut_mask = 16'hAACC;
defparam \td_shift~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~16 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~15_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~16_combout ),
	.cout());
defparam \td_shift~16 .lut_mask = 16'hACFF;
defparam \td_shift~16 .sum_lutc_input = "datac";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~16_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cycloneive_lcell_comb \td_shift~13 (
	.dataa(\td_shift[5]~q ),
	.datab(\rdata[2]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~13_combout ),
	.cout());
defparam \td_shift~13 .lut_mask = 16'hACAC;
defparam \td_shift~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~14 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~1_combout ),
	.datad(\td_shift~13_combout ),
	.cin(gnd),
	.combout(\td_shift~14_combout ),
	.cout());
defparam \td_shift~14 .lut_mask = 16'hFFEF;
defparam \td_shift~14 .sum_lutc_input = "datac";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~14_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cycloneive_lcell_comb \td_shift~11 (
	.dataa(\td_shift[4]~q ),
	.datab(\rdata[1]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~11_combout ),
	.cout());
defparam \td_shift~11 .lut_mask = 16'hACAC;
defparam \td_shift~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~12 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~1_combout ),
	.datad(\td_shift~11_combout ),
	.cin(gnd),
	.combout(\td_shift~12_combout ),
	.cout());
defparam \td_shift~12 .lut_mask = 16'hFFEF;
defparam \td_shift~12 .sum_lutc_input = "datac";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~12_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

cycloneive_lcell_comb \td_shift~8 (
	.dataa(\td_shift[3]~q ),
	.datab(\rdata[0]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~8_combout ),
	.cout());
defparam \td_shift~8 .lut_mask = 16'hAACC;
defparam \td_shift~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~9 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~8_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~9_combout ),
	.cout());
defparam \td_shift~9 .lut_mask = 16'hACFF;
defparam \td_shift~9 .sum_lutc_input = "datac";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cycloneive_lcell_comb \write_stalled~2 (
	.dataa(\write_stalled~q ),
	.datab(\td_shift[10]~q ),
	.datac(altera_internal_jtag1),
	.datad(\tck_t_dav~q ),
	.cin(gnd),
	.combout(\write_stalled~2_combout ),
	.cout());
defparam \write_stalled~2 .lut_mask = 16'hEFFF;
defparam \write_stalled~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_stalled~4 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(virtual_ir_scan_reg),
	.datac(irf_reg_0_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_stalled~4_combout ),
	.cout());
defparam \write_stalled~4 .lut_mask = 16'hBFBF;
defparam \write_stalled~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_stalled~3 (
	.dataa(\count[1]~q ),
	.datab(\state~q ),
	.datac(state_4),
	.datad(\write_stalled~4_combout ),
	.cin(gnd),
	.combout(\write_stalled~3_combout ),
	.cout());
defparam \write_stalled~3 .lut_mask = 16'hFFFE;
defparam \write_stalled~3 .sum_lutc_input = "datac";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cycloneive_lcell_comb \td_shift~5 (
	.dataa(\td_shift[2]~q ),
	.datab(\write_stalled~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~5_combout ),
	.cout());
defparam \td_shift~5 .lut_mask = 16'hAACC;
defparam \td_shift~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~6 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~5_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~6_combout ),
	.cout());
defparam \td_shift~6 .lut_mask = 16'hACFF;
defparam \td_shift~6 .sum_lutc_input = "datac";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cycloneive_lcell_comb \td_shift~0 (
	.dataa(\td_shift[1]~q ),
	.datab(\rvalid~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~0_combout ),
	.cout());
defparam \td_shift~0 .lut_mask = 16'hAACC;
defparam \td_shift~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~2 (
	.dataa(\td_shift~1_combout ),
	.datab(altera_internal_jtag1),
	.datac(\state~q ),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\td_shift~2_combout ),
	.cout());
defparam \td_shift~2 .lut_mask = 16'hEFFF;
defparam \td_shift~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~3 (
	.dataa(\tck_t_dav~q ),
	.datab(\td_shift~0_combout ),
	.datac(\td_shift~2_combout ),
	.datad(\state~q ),
	.cin(gnd),
	.combout(\td_shift~3_combout ),
	.cout());
defparam \td_shift~3 .lut_mask = 16'hACFF;
defparam \td_shift~3 .sum_lutc_input = "datac";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cycloneive_lcell_comb \rvalid0~0 (
	.dataa(rvalid01),
	.datab(r_val),
	.datac(r_ena11),
	.datad(gnd),
	.cin(gnd),
	.combout(\rvalid0~0_combout ),
	.cout());
defparam \rvalid0~0 .lut_mask = 16'h7F7F;
defparam \rvalid0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h5555;
defparam \read~0 .sum_lutc_input = "datac";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cycloneive_lcell_comb \rvalid0~1 (
	.dataa(\read1~q ),
	.datab(\read2~q ),
	.datac(\user_saw_rvalid~q ),
	.datad(\read_req~q ),
	.cin(gnd),
	.combout(\rvalid0~1_combout ),
	.cout());
defparam \rvalid0~1 .lut_mask = 16'h6FFF;
defparam \rvalid0~1 .sum_lutc_input = "datac";

dffeas rst2(
	.clk(clk),
	.d(rst11),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cycloneive_lcell_comb \rvalid0~2 (
	.dataa(\rvalid0~0_combout ),
	.datab(\rvalid0~1_combout ),
	.datac(gnd),
	.datad(\rst2~q ),
	.cin(gnd),
	.combout(\rvalid0~2_combout ),
	.cout());
defparam \rvalid0~2 .lut_mask = 16'hDDFF;
defparam \rvalid0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~4 (
	.dataa(\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\write~4_combout ),
	.cout());
defparam \write~4 .lut_mask = 16'h5555;
defparam \write~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~3 (
	.dataa(\count[8]~q ),
	.datab(\state~q ),
	.datac(state_4),
	.datad(\write_stalled~4_combout ),
	.cin(gnd),
	.combout(\write~3_combout ),
	.cout());
defparam \write~3 .lut_mask = 16'hFFFE;
defparam \write~3 .sum_lutc_input = "datac";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~4_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~3_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cycloneive_lcell_comb \t_ena~2 (
	.dataa(t_ena1),
	.datab(\write_valid~q ),
	.datac(t_dav),
	.datad(\write_stalled~q ),
	.cin(gnd),
	.combout(\t_ena~2_combout ),
	.cout());
defparam \t_ena~2 .lut_mask = 16'hEFFF;
defparam \t_ena~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \t_ena~3 (
	.dataa(\write1~q ),
	.datab(\write2~q ),
	.datac(\rst2~q ),
	.datad(\t_ena~2_combout ),
	.cin(gnd),
	.combout(\t_ena~3_combout ),
	.cout());
defparam \t_ena~3 .lut_mask = 16'hFFF6;
defparam \t_ena~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\write1~q ),
	.datad(\write2~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'h0FF0;
defparam \always2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \t_pause~0 (
	.dataa(\always2~0_combout ),
	.datab(t_dav),
	.datac(\write_stalled~q ),
	.datad(\write_valid~q ),
	.cin(gnd),
	.combout(\t_pause~0_combout ),
	.cout());
defparam \t_pause~0 .lut_mask = 16'hFEFF;
defparam \t_pause~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jupdate~0 (
	.dataa(\jupdate~q ),
	.datab(irf_reg_0_1),
	.datac(\always0~0_combout ),
	.datad(state_8),
	.cin(gnd),
	.combout(\jupdate~0_combout ),
	.cout());
defparam \jupdate~0 .lut_mask = 16'h6996;
defparam \jupdate~0 .sum_lutc_input = "datac";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cycloneive_lcell_comb \t_pause~1 (
	.dataa(\rst2~q ),
	.datab(\t_pause~0_combout ),
	.datac(\jupdate1~q ),
	.datad(\jupdate2~q ),
	.cin(gnd),
	.combout(\t_pause~1_combout ),
	.cout());
defparam \t_pause~1 .lut_mask = 16'hEFFE;
defparam \t_pause~1 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_jtag_scfifo_r (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	altera_reset_synchronizer_int_chain_out,
	b_full,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wr_rfifo,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wr_rfifo;
input 	wdata_0;
input 	wdata_1;
input 	wdata_2;
input 	wdata_3;
input 	wdata_4;
input 	wdata_5;
input 	wdata_6;
input 	wdata_7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_1 rfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wrreq(wr_rfifo),
	.data({wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.clock(clk_clk));

endmodule

module niosII_scfifo_1 (
	q,
	altera_reset_synchronizer_int_chain_out,
	b_full,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_jr21 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module niosII_scfifo_jr21 (
	q,
	altera_reset_synchronizer_int_chain_out,
	b_full,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_a_dpfifo_l011 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module niosII_a_dpfifo_l011 (
	q,
	altera_reset_synchronizer_int_chain_out,
	b_full,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


niosII_a_fefifo_7cf fifo_state(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_full1(b_full),
	.b_non_empty1(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wreq(wreq),
	.clock(clock));

niosII_cntr_1ob_1 wr_ptr(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

niosII_cntr_1ob rd_ptr_count(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.fifo_rd(fifo_rd),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

niosII_altsyncram_nio1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(fifo_rd),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

endmodule

module niosII_a_fefifo_7cf (
	altera_reset_synchronizer_int_chain_out,
	b_full1,
	b_non_empty1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wreq,
	clock)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_full1;
output 	b_non_empty1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~4_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;
wire \b_non_empty~0_combout ;
wire \_~2_combout ;
wire \_~3_combout ;
wire \b_non_empty~1_combout ;


niosII_cntr_do7 count_usedw(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.updown(wreq),
	._(\_~4_combout ),
	.clock(clock));

cycloneive_lcell_comb \_~4 (
	.dataa(t_ena),
	.datab(b_full1),
	.datac(fifo_rd),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'h9696;
defparam \_~4 .sum_lutc_input = "datac";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cycloneive_lcell_comb \b_full~0 (
	.dataa(b_non_empty1),
	.datab(counter_reg_bit_5),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_3),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_0),
	.datad(t_ena),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(fifo_rd),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~0 (
	.dataa(b_full1),
	.datab(t_ena),
	.datac(gnd),
	.datad(b_non_empty1),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hEEFF;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_5),
	.datab(counter_reg_bit_4),
	.datac(wreq),
	.datad(fifo_rd),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hFEFF;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~1 (
	.dataa(\b_non_empty~0_combout ),
	.datab(b_non_empty1),
	.datac(\_~2_combout ),
	.datad(\_~3_combout ),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hFFFE;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

endmodule

module niosII_cntr_do7 (
	altera_reset_synchronizer_int_chain_out,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	updown,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	updown;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_altsyncram_nio1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_r:the_niosII_jtag_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_r:the_niosII_jtag_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_r:the_niosII_jtag_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_r:the_niosII_jtag_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_r:the_niosII_jtag_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_r:the_niosII_jtag_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_r:the_niosII_jtag_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_r:the_niosII_jtag_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module niosII_cntr_1ob (
	altera_reset_synchronizer_int_chain_out,
	fifo_rd,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
input 	fifo_rd;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_cntr_1ob_1 (
	altera_reset_synchronizer_int_chain_out,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_niosII_jtag_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	altera_reset_synchronizer_int_chain_out,
	b_non_empty,
	r_val,
	fifo_wr,
	out_data_buffer_7,
	out_data_buffer_0,
	b_full,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_non_empty;
input 	r_val;
input 	fifo_wr;
input 	out_data_buffer_7;
input 	out_data_buffer_0;
output 	b_full;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
input 	out_data_buffer_1;
input 	out_data_buffer_2;
input 	out_data_buffer_3;
input 	out_data_buffer_4;
input 	out_data_buffer_5;
input 	out_data_buffer_6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_2 wfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(fifo_wr),
	.data({out_data_buffer_7,out_data_buffer_6,out_data_buffer_5,out_data_buffer_4,out_data_buffer_3,out_data_buffer_2,out_data_buffer_1,out_data_buffer_0}),
	.b_full(b_full),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.clock(clk_clk));

endmodule

module niosII_scfifo_2 (
	q,
	altera_reset_synchronizer_int_chain_out,
	b_non_empty,
	r_val,
	wrreq,
	data,
	b_full,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_0,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
input 	[7:0] data;
output 	b_full;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_jr21_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.b_full(b_full),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.clock(clock));

endmodule

module niosII_scfifo_jr21_1 (
	q,
	altera_reset_synchronizer_int_chain_out,
	b_non_empty,
	r_val,
	wrreq,
	data,
	b_full,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_0,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
input 	[7:0] data;
output 	b_full;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_a_dpfifo_l011_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.b_full(b_full),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.clock(clock));

endmodule

module niosII_a_dpfifo_l011_1 (
	q,
	altera_reset_synchronizer_int_chain_out,
	b_non_empty,
	r_val,
	wreq,
	data,
	b_full,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_0,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_non_empty;
input 	r_val;
input 	wreq;
input 	[7:0] data;
output 	b_full;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


niosII_cntr_1ob_3 wr_ptr(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

niosII_cntr_1ob_2 rd_ptr_count(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.r_val(r_val),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

niosII_altsyncram_nio1_1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(r_val),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

niosII_a_fefifo_7cf_1 fifo_state(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.b_non_empty1(b_non_empty),
	.r_val(r_val),
	.wreq(wreq),
	.b_full1(b_full),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.clock(clock));

endmodule

module niosII_a_fefifo_7cf_1 (
	altera_reset_synchronizer_int_chain_out,
	b_non_empty1,
	r_val,
	wreq,
	b_full1,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	b_non_empty1;
input 	r_val;
input 	wreq;
output 	b_full1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;


niosII_cntr_do7_1 count_usedw(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.updown(wreq),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	._(\_~0_combout ),
	.clock(clock));

cycloneive_lcell_comb \_~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(wreq),
	.datad(r_val),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h0FF0;
defparam \_~0 .sum_lutc_input = "datac";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

cycloneive_lcell_comb \b_non_empty~0 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hFFFE;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~1 (
	.dataa(\b_non_empty~0_combout ),
	.datab(counter_reg_bit_3),
	.datac(r_val),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hEFFF;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~2 (
	.dataa(wreq),
	.datab(b_full1),
	.datac(b_non_empty1),
	.datad(\b_non_empty~1_combout ),
	.cin(gnd),
	.combout(\b_non_empty~2_combout ),
	.cout());
defparam \b_non_empty~2 .lut_mask = 16'hFFFE;
defparam \b_non_empty~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~0 (
	.dataa(wreq),
	.datab(b_non_empty1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(r_val),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

endmodule

module niosII_cntr_do7_1 (
	altera_reset_synchronizer_int_chain_out,
	updown,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_0,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
input 	updown;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_altsyncram_nio1_1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_w:the_niosII_jtag_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_w:the_niosII_jtag_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_w:the_niosII_jtag_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_w:the_niosII_jtag_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_w:the_niosII_jtag_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_w:the_niosII_jtag_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_w:the_niosII_jtag_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosII_jtag:jtag|niosII_jtag_scfifo_w:the_niosII_jtag_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

endmodule

module niosII_cntr_1ob_2 (
	altera_reset_synchronizer_int_chain_out,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_cntr_1ob_3 (
	altera_reset_synchronizer_int_chain_out,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_niosII_mm_interconnect_0 (
	wire_pll7_clk_0,
	W_alu_result_6,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_5,
	W_alu_result_7,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	byteen_reg_0,
	byteen_reg_1,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	readdata_0,
	readdata_01,
	readdata_4,
	readdata_1,
	readdata_11,
	readdata_23,
	readdata_231,
	readdata_22,
	readdata_221,
	readdata_21,
	readdata_211,
	readdata_20,
	readdata_201,
	readdata_19,
	readdata_191,
	readdata_18,
	readdata_181,
	readdata_17,
	readdata_171,
	readdata_16,
	readdata_161,
	r_sync_rst,
	r_sync_rst1,
	saved_grant_0,
	saved_grant_1,
	out_data_buffer_38,
	src_data_38,
	src_data_39,
	src_data_40,
	src_payload,
	entries_1,
	entries_0,
	mem_used_1,
	d_read,
	read_accepted,
	hold_waitrequest,
	d_write,
	write_accepted,
	cp_valid,
	Equal3,
	m0_read,
	m0_write,
	src_payload1,
	mem_used_11,
	wait_latency_counter_1,
	src_valid,
	src_valid1,
	src_data_46,
	out_data_buffer_65,
	p1_wr_strobe,
	src_payload2,
	d_writedata_0,
	d_byteenable_0,
	Equal9,
	read_latency_shift_reg,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	out_data_buffer_0,
	out_data_toggle_flopped,
	dreg_0,
	mem_used_12,
	wire_pfdena_reg_ena,
	out_data_buffer_651,
	out_data_buffer_381,
	out_data_buffer_39,
	altera_reset_synchronizer_int_chain_out,
	saved_grant_01,
	d_byteenable_1,
	use_reg,
	saved_grant_11,
	WideOr0,
	Equal0,
	i_read,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	Equal1,
	Equal4,
	WideOr1,
	m0_write1,
	mem_used_7,
	src_data_66,
	F_pc_8,
	out_data_28,
	src_valid2,
	src12_valid,
	m0_write2,
	out_data_42,
	F_pc_9,
	out_data_29,
	out_data_31,
	out_data_30,
	out_data_33,
	out_data_32,
	out_data_35,
	out_data_34,
	out_data_37,
	out_data_36,
	out_data_39,
	out_data_38,
	out_data_41,
	out_data_40,
	out_data_19,
	F_pc_0,
	out_data_20,
	F_pc_1,
	out_data_21,
	F_pc_2,
	out_data_22,
	F_pc_3,
	out_data_23,
	F_pc_4,
	out_data_24,
	F_pc_5,
	out_data_25,
	F_pc_6,
	out_data_26,
	F_pc_7,
	out_data_27,
	always0,
	waitrequest,
	mem_84_0,
	mem_66_0,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	mem_54_0,
	src0_valid,
	WideOr11,
	mem_used_13,
	wait_latency_counter_0,
	wait_latency_counter_11,
	read_latency_shift_reg1,
	write,
	Equal12,
	mem_used_14,
	saved_grant_02,
	waitrequest1,
	mem_used_15,
	cpu_data_master_waitrequest,
	src_payload3,
	src_data_661,
	av_begintransfer,
	d_writedata_10,
	src_payload4,
	rst1,
	out_data_buffer_66,
	d_byteenable_2,
	d_byteenable_3,
	src1_valid,
	read_accepted1,
	src1_valid1,
	hbreak_enabled,
	read_latency_shift_reg2,
	d_writedata_8,
	d_writedata_9,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	WideOr12,
	write1,
	Equal121,
	rf_source_valid,
	uav_write,
	src_payload5,
	out_valid,
	av_readdata_pre_0,
	out_data_buffer_01,
	data_reg_0,
	out_payload_0,
	source_addr_1,
	F_iw_0,
	av_readdata_pre_1,
	out_data_buffer_1,
	out_payload_1,
	src_data_1,
	av_readdata_pre_2,
	out_data_buffer_2,
	data_reg_2,
	out_payload_2,
	F_iw_2,
	av_readdata_pre_3,
	out_data_buffer_3,
	out_payload_3,
	src_data_3,
	av_readdata_pre_4,
	out_data_buffer_4,
	out_payload_4,
	src_data_4,
	read_latency_shift_reg3,
	b_full,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	period_l_wr_strobe,
	src_data_461,
	out_data_toggle_flopped1,
	av_readdata_pre_11,
	out_data_buffer_11,
	out_payload_11,
	src_data_11,
	av_readdata_pre_13,
	out_data_buffer_13,
	out_payload_13,
	src_data_13,
	av_readdata_pre_16,
	out_data_buffer_16,
	src_payload6,
	av_readdata_pre_12,
	out_data_buffer_12,
	data_reg_12,
	out_payload_12,
	F_iw_12,
	av_readdata_pre_5,
	out_data_buffer_5,
	out_payload_5,
	src_data_5,
	av_readdata_pre_14,
	out_data_buffer_14,
	data_reg_14,
	out_payload_14,
	F_iw_14,
	av_readdata_pre_15,
	out_data_buffer_15,
	out_payload_15,
	src_data_15,
	av_readdata_pre_10,
	out_data_buffer_10,
	data_reg_10,
	out_payload_10,
	F_iw_10,
	av_readdata_pre_9,
	out_data_buffer_9,
	data_reg_9,
	out_payload_9,
	F_iw_9,
	av_readdata_pre_8,
	out_data_buffer_8,
	data_reg_8,
	out_payload_8,
	F_iw_8,
	av_readdata_pre_7,
	out_data_buffer_7,
	data_reg_7,
	out_payload_7,
	F_iw_7,
	av_readdata_pre_6,
	out_data_buffer_6,
	data_reg_6,
	out_payload_6,
	F_iw_6,
	av_readdata_pre_21,
	out_data_buffer_21,
	av_readdata_pre_30,
	out_data_buffer_30,
	av_readdata_pre_29,
	out_data_buffer_29,
	av_readdata_pre_28,
	out_data_buffer_28,
	av_readdata_pre_27,
	out_data_buffer_27,
	av_readdata_pre_26,
	out_data_buffer_26,
	av_readdata_pre_25,
	out_data_buffer_25,
	av_readdata_pre_24,
	out_data_buffer_24,
	av_readdata_pre_23,
	out_data_buffer_23,
	av_readdata_pre_22,
	out_data_buffer_22,
	av_readdata_pre_20,
	out_data_buffer_20,
	av_readdata_pre_19,
	out_data_buffer_19,
	av_readdata_pre_18,
	out_data_buffer_18,
	av_readdata_pre_17,
	out_data_buffer_17,
	src_payload7,
	readdata_02,
	readdata_03,
	readdata_04,
	readdata_05,
	out_valid1,
	src_data_0,
	readdata_06,
	readdata_12,
	readdata_2,
	readdata_3,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_110,
	src_data_12,
	src_data_2,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_27,
	readdata_28,
	src_data_21,
	readdata_31,
	readdata_32,
	readdata_33,
	readdata_34,
	readdata_35,
	src_data_31,
	readdata_41,
	readdata_42,
	readdata_43,
	readdata_44,
	av_readdata_pre_301,
	src_data_41,
	readdata_5,
	readdata_51,
	readdata_52,
	readdata_53,
	src_data_51,
	readdata_6,
	readdata_61,
	readdata_62,
	readdata_63,
	src_data_6,
	readdata_7,
	readdata_71,
	readdata_72,
	readdata_73,
	src_data_7,
	src_payload8,
	src_payload9,
	src_data_381,
	src_data_391,
	src_data_401,
	src_data_411,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	dreg_01,
	av_waitrequest,
	mem_used_16,
	out_data_buffer_661,
	out_data_buffer_382,
	out_data_buffer_71,
	za_valid,
	readdata_111,
	readdata_131,
	readdata_162,
	readdata_121,
	readdata_54,
	readdata_141,
	readdata_151,
	readdata_10,
	av_readdata_pre_31,
	out_data_buffer_31,
	readdata_9,
	readdata_8,
	readdata_74,
	readdata_64,
	out_data_buffer_261,
	readdata_212,
	readdata_30,
	out_data_buffer_251,
	src_payload10,
	readdata_29,
	out_data_buffer_241,
	readdata_281,
	readdata_232,
	src_payload11,
	readdata_271,
	readdata_222,
	src_payload12,
	readdata_261,
	readdata_213,
	src_payload13,
	readdata_251,
	readdata_202,
	src_payload14,
	readdata_241,
	readdata_192,
	src_payload15,
	readdata_233,
	readdata_182,
	src_payload16,
	readdata_223,
	readdata_172,
	src_payload17,
	readdata_163,
	src_payload18,
	readdata_203,
	readdata_152,
	readdata_153,
	readdata_154,
	src_data_151,
	readdata_193,
	readdata_142,
	src_data_14,
	readdata_183,
	readdata_132,
	src_data_131,
	readdata_173,
	readdata_122,
	src_data_121,
	readdata_112,
	src_data_111,
	readdata_101,
	src_data_10,
	readdata_91,
	readdata_92,
	readdata_93,
	src_data_9,
	readdata_81,
	readdata_82,
	readdata_83,
	src_data_8,
	src_payload19,
	av_readdata_pre_01,
	readdata_07,
	readdata_08,
	readdata_113,
	readdata_114,
	readdata_210,
	readdata_214,
	readdata_36,
	readdata_37,
	readdata_45,
	readdata_46,
	readdata_55,
	readdata_56,
	readdata_65,
	readdata_66,
	readdata_75,
	readdata_76,
	src_payload20,
	out_data_buffer_652,
	out_data_buffer_02,
	b_full1,
	counter_reg_bit_21,
	counter_reg_bit_11,
	counter_reg_bit_51,
	counter_reg_bit_41,
	counter_reg_bit_31,
	counter_reg_bit_01,
	out_data_buffer_271,
	out_data_buffer_281,
	out_data_buffer_291,
	out_data_buffer_301,
	out_data_buffer_311,
	readdata_311,
	readdata_155,
	readdata_156,
	readdata_143,
	readdata_133,
	readdata_123,
	readdata_115,
	readdata_116,
	readdata_102,
	readdata_103,
	readdata_94,
	readdata_95,
	readdata_84,
	readdata_85,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	readdata_09,
	za_data_0,
	readdata_117,
	za_data_1,
	readdata_215,
	za_data_2,
	readdata_38,
	za_data_3,
	readdata_47,
	za_data_4,
	out_data_buffer_110,
	readdata_118,
	za_data_11,
	readdata_134,
	za_data_13,
	readdata_164,
	readdata_124,
	za_data_12,
	readdata_57,
	za_data_5,
	readdata_144,
	za_data_14,
	readdata_157,
	za_data_15,
	readdata_104,
	za_data_10,
	readdata_96,
	za_data_9,
	readdata_86,
	za_data_8,
	readdata_77,
	za_data_7,
	readdata_67,
	za_data_6,
	readdata_216,
	readdata_301,
	readdata_291,
	readdata_282,
	readdata_272,
	readdata_262,
	readdata_252,
	readdata_242,
	readdata_234,
	readdata_224,
	readdata_204,
	readdata_194,
	readdata_184,
	readdata_174,
	src_payload25,
	read_0,
	av_readdata_0,
	readdata_010,
	av_readdata_9,
	src_data_412,
	src_data_421,
	src_data_431,
	src_data_441,
	src_data_451,
	src_payload26,
	av_readdata_1,
	readdata_119,
	av_readdata_2,
	av_readdata_3,
	av_readdata_4,
	av_readdata_5,
	av_readdata_6,
	av_readdata_7,
	out_data_buffer_210,
	src_payload27,
	src_data_33,
	src_payload28,
	src_payload29,
	src_data_34,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	readdata_312,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_data_35,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_payload46,
	src_payload47,
	src_payload48,
	src_payload49,
	rvalid,
	src_payload50,
	woverflow,
	src_payload51,
	src_payload52,
	ac,
	av_readdata_8,
	out_data_buffer_111,
	out_data_buffer_32,
	src_payload53,
	src_payload54,
	src_payload55,
	src_payload56,
	src_payload57,
	src_payload58,
	src_payload59,
	src_payload60,
	out_data_buffer_101,
	out_data_buffer_41,
	out_data_buffer_51,
	out_data_buffer_61,
	write2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_6;
input 	W_alu_result_26;
input 	W_alu_result_25;
input 	W_alu_result_24;
input 	W_alu_result_23;
input 	W_alu_result_22;
input 	W_alu_result_21;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_5;
input 	W_alu_result_7;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
output 	byteen_reg_0;
output 	byteen_reg_1;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	readdata_0;
input 	readdata_01;
input 	readdata_4;
input 	readdata_1;
input 	readdata_11;
input 	readdata_23;
input 	readdata_231;
input 	readdata_22;
input 	readdata_221;
input 	readdata_21;
input 	readdata_211;
input 	readdata_20;
input 	readdata_201;
input 	readdata_19;
input 	readdata_191;
input 	readdata_18;
input 	readdata_181;
input 	readdata_17;
input 	readdata_171;
input 	readdata_16;
input 	readdata_161;
input 	r_sync_rst;
input 	r_sync_rst1;
output 	saved_grant_0;
output 	saved_grant_1;
output 	out_data_buffer_38;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_payload;
input 	entries_1;
input 	entries_0;
output 	mem_used_1;
input 	d_read;
output 	read_accepted;
output 	hold_waitrequest;
input 	d_write;
output 	write_accepted;
output 	cp_valid;
output 	Equal3;
output 	m0_read;
output 	m0_write;
output 	src_payload1;
output 	mem_used_11;
output 	wait_latency_counter_1;
output 	src_valid;
output 	src_valid1;
output 	src_data_46;
output 	out_data_buffer_65;
input 	p1_wr_strobe;
output 	src_payload2;
input 	d_writedata_0;
input 	d_byteenable_0;
output 	Equal9;
output 	read_latency_shift_reg;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	out_data_buffer_0;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	mem_used_12;
input 	wire_pfdena_reg_ena;
output 	out_data_buffer_651;
output 	out_data_buffer_381;
output 	out_data_buffer_39;
input 	altera_reset_synchronizer_int_chain_out;
output 	saved_grant_01;
input 	d_byteenable_1;
output 	use_reg;
output 	saved_grant_11;
output 	WideOr0;
input 	Equal0;
input 	i_read;
input 	F_pc_24;
input 	F_pc_23;
input 	F_pc_22;
input 	F_pc_21;
input 	F_pc_20;
input 	F_pc_19;
input 	F_pc_18;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
input 	F_pc_10;
output 	Equal1;
output 	Equal4;
output 	WideOr1;
output 	m0_write1;
output 	mem_used_7;
output 	src_data_66;
input 	F_pc_8;
output 	out_data_28;
output 	src_valid2;
output 	src12_valid;
output 	m0_write2;
output 	out_data_42;
input 	F_pc_9;
output 	out_data_29;
output 	out_data_31;
output 	out_data_30;
output 	out_data_33;
output 	out_data_32;
output 	out_data_35;
output 	out_data_34;
output 	out_data_37;
output 	out_data_36;
output 	out_data_39;
output 	out_data_38;
output 	out_data_41;
output 	out_data_40;
output 	out_data_19;
input 	F_pc_0;
output 	out_data_20;
input 	F_pc_1;
output 	out_data_21;
input 	F_pc_2;
output 	out_data_22;
input 	F_pc_3;
output 	out_data_23;
input 	F_pc_4;
output 	out_data_24;
input 	F_pc_5;
output 	out_data_25;
input 	F_pc_6;
output 	out_data_26;
input 	F_pc_7;
output 	out_data_27;
input 	always0;
input 	waitrequest;
output 	mem_84_0;
output 	mem_66_0;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg_01;
output 	read_latency_shift_reg_02;
output 	mem_54_0;
output 	src0_valid;
output 	WideOr11;
output 	mem_used_13;
output 	wait_latency_counter_0;
output 	wait_latency_counter_11;
output 	read_latency_shift_reg1;
output 	write;
output 	Equal12;
output 	mem_used_14;
output 	saved_grant_02;
input 	waitrequest1;
output 	mem_used_15;
output 	cpu_data_master_waitrequest;
output 	src_payload3;
output 	src_data_661;
output 	av_begintransfer;
input 	d_writedata_10;
output 	src_payload4;
input 	rst1;
output 	out_data_buffer_66;
input 	d_byteenable_2;
input 	d_byteenable_3;
output 	src1_valid;
output 	read_accepted1;
output 	src1_valid1;
input 	hbreak_enabled;
output 	read_latency_shift_reg2;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
output 	WideOr12;
output 	write1;
output 	Equal121;
output 	rf_source_valid;
output 	uav_write;
output 	src_payload5;
output 	out_valid;
output 	av_readdata_pre_0;
output 	out_data_buffer_01;
output 	data_reg_0;
output 	out_payload_0;
output 	source_addr_1;
input 	F_iw_0;
output 	av_readdata_pre_1;
output 	out_data_buffer_1;
output 	out_payload_1;
output 	src_data_1;
output 	av_readdata_pre_2;
output 	out_data_buffer_2;
output 	data_reg_2;
output 	out_payload_2;
input 	F_iw_2;
output 	av_readdata_pre_3;
output 	out_data_buffer_3;
output 	out_payload_3;
output 	src_data_3;
output 	av_readdata_pre_4;
output 	out_data_buffer_4;
output 	out_payload_4;
output 	src_data_4;
output 	read_latency_shift_reg3;
input 	b_full;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
input 	period_l_wr_strobe;
output 	src_data_461;
output 	out_data_toggle_flopped1;
output 	av_readdata_pre_11;
output 	out_data_buffer_11;
output 	out_payload_11;
output 	src_data_11;
output 	av_readdata_pre_13;
output 	out_data_buffer_13;
output 	out_payload_13;
output 	src_data_13;
output 	av_readdata_pre_16;
output 	out_data_buffer_16;
output 	src_payload6;
output 	av_readdata_pre_12;
output 	out_data_buffer_12;
output 	data_reg_12;
output 	out_payload_12;
input 	F_iw_12;
output 	av_readdata_pre_5;
output 	out_data_buffer_5;
output 	out_payload_5;
output 	src_data_5;
output 	av_readdata_pre_14;
output 	out_data_buffer_14;
output 	data_reg_14;
output 	out_payload_14;
input 	F_iw_14;
output 	av_readdata_pre_15;
output 	out_data_buffer_15;
output 	out_payload_15;
output 	src_data_15;
output 	av_readdata_pre_10;
output 	out_data_buffer_10;
output 	data_reg_10;
output 	out_payload_10;
input 	F_iw_10;
output 	av_readdata_pre_9;
output 	out_data_buffer_9;
output 	data_reg_9;
output 	out_payload_9;
input 	F_iw_9;
output 	av_readdata_pre_8;
output 	out_data_buffer_8;
output 	data_reg_8;
output 	out_payload_8;
input 	F_iw_8;
output 	av_readdata_pre_7;
output 	out_data_buffer_7;
output 	data_reg_7;
output 	out_payload_7;
input 	F_iw_7;
output 	av_readdata_pre_6;
output 	out_data_buffer_6;
output 	data_reg_6;
output 	out_payload_6;
input 	F_iw_6;
output 	av_readdata_pre_21;
output 	out_data_buffer_21;
output 	av_readdata_pre_30;
output 	out_data_buffer_30;
output 	av_readdata_pre_29;
output 	out_data_buffer_29;
output 	av_readdata_pre_28;
output 	out_data_buffer_28;
output 	av_readdata_pre_27;
output 	out_data_buffer_27;
output 	av_readdata_pre_26;
output 	out_data_buffer_26;
output 	av_readdata_pre_25;
output 	out_data_buffer_25;
output 	av_readdata_pre_24;
output 	out_data_buffer_24;
output 	av_readdata_pre_23;
output 	out_data_buffer_23;
output 	av_readdata_pre_22;
output 	out_data_buffer_22;
output 	av_readdata_pre_20;
output 	out_data_buffer_20;
output 	av_readdata_pre_19;
output 	out_data_buffer_19;
output 	av_readdata_pre_18;
output 	out_data_buffer_18;
output 	av_readdata_pre_17;
output 	out_data_buffer_17;
output 	src_payload7;
input 	readdata_02;
input 	readdata_03;
input 	readdata_04;
input 	readdata_05;
output 	out_valid1;
output 	src_data_0;
input 	readdata_06;
input 	readdata_12;
input 	readdata_2;
input 	readdata_3;
input 	readdata_13;
input 	readdata_14;
input 	readdata_15;
input 	readdata_110;
output 	src_data_12;
output 	src_data_2;
input 	readdata_24;
input 	readdata_25;
input 	readdata_26;
input 	readdata_27;
input 	readdata_28;
output 	src_data_21;
input 	readdata_31;
input 	readdata_32;
input 	readdata_33;
input 	readdata_34;
input 	readdata_35;
output 	src_data_31;
input 	readdata_41;
input 	readdata_42;
input 	readdata_43;
input 	readdata_44;
output 	av_readdata_pre_301;
output 	src_data_41;
input 	readdata_5;
input 	readdata_51;
input 	readdata_52;
input 	readdata_53;
output 	src_data_51;
input 	readdata_6;
input 	readdata_61;
input 	readdata_62;
input 	readdata_63;
output 	src_data_6;
input 	readdata_7;
input 	readdata_71;
input 	readdata_72;
input 	readdata_73;
output 	src_data_7;
output 	src_payload8;
output 	src_payload9;
output 	src_data_381;
output 	src_data_391;
output 	src_data_401;
output 	src_data_411;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_32;
input 	b_non_empty;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
output 	dreg_01;
input 	av_waitrequest;
output 	mem_used_16;
output 	out_data_buffer_661;
output 	out_data_buffer_382;
output 	out_data_buffer_71;
input 	za_valid;
input 	readdata_111;
input 	readdata_131;
input 	readdata_162;
input 	readdata_121;
input 	readdata_54;
input 	readdata_141;
input 	readdata_151;
input 	readdata_10;
output 	av_readdata_pre_31;
output 	out_data_buffer_31;
input 	readdata_9;
input 	readdata_8;
input 	readdata_74;
input 	readdata_64;
output 	out_data_buffer_261;
input 	readdata_212;
input 	readdata_30;
output 	out_data_buffer_251;
output 	src_payload10;
input 	readdata_29;
output 	out_data_buffer_241;
input 	readdata_281;
input 	readdata_232;
output 	src_payload11;
input 	readdata_271;
input 	readdata_222;
output 	src_payload12;
input 	readdata_261;
input 	readdata_213;
output 	src_payload13;
input 	readdata_251;
input 	readdata_202;
output 	src_payload14;
input 	readdata_241;
input 	readdata_192;
output 	src_payload15;
input 	readdata_233;
input 	readdata_182;
output 	src_payload16;
input 	readdata_223;
input 	readdata_172;
output 	src_payload17;
input 	readdata_163;
output 	src_payload18;
input 	readdata_203;
input 	readdata_152;
input 	readdata_153;
input 	readdata_154;
output 	src_data_151;
input 	readdata_193;
input 	readdata_142;
output 	src_data_14;
input 	readdata_183;
input 	readdata_132;
output 	src_data_131;
input 	readdata_173;
input 	readdata_122;
output 	src_data_121;
input 	readdata_112;
output 	src_data_111;
input 	readdata_101;
output 	src_data_10;
input 	readdata_91;
input 	readdata_92;
input 	readdata_93;
output 	src_data_9;
input 	readdata_81;
input 	readdata_82;
input 	readdata_83;
output 	src_data_8;
output 	src_payload19;
output 	av_readdata_pre_01;
input 	readdata_07;
input 	readdata_08;
input 	readdata_113;
input 	readdata_114;
input 	readdata_210;
input 	readdata_214;
input 	readdata_36;
input 	readdata_37;
input 	readdata_45;
input 	readdata_46;
input 	readdata_55;
input 	readdata_56;
input 	readdata_65;
input 	readdata_66;
input 	readdata_75;
input 	readdata_76;
output 	src_payload20;
output 	out_data_buffer_652;
output 	out_data_buffer_02;
input 	b_full1;
input 	counter_reg_bit_21;
input 	counter_reg_bit_11;
input 	counter_reg_bit_51;
input 	counter_reg_bit_41;
input 	counter_reg_bit_31;
input 	counter_reg_bit_01;
output 	out_data_buffer_271;
output 	out_data_buffer_281;
output 	out_data_buffer_291;
output 	out_data_buffer_301;
output 	out_data_buffer_311;
input 	readdata_311;
input 	readdata_155;
input 	readdata_156;
input 	readdata_143;
input 	readdata_133;
input 	readdata_123;
input 	readdata_115;
input 	readdata_116;
input 	readdata_102;
input 	readdata_103;
input 	readdata_94;
input 	readdata_95;
input 	readdata_84;
input 	readdata_85;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
input 	readdata_09;
input 	za_data_0;
input 	readdata_117;
input 	za_data_1;
input 	readdata_215;
input 	za_data_2;
input 	readdata_38;
input 	za_data_3;
input 	readdata_47;
input 	za_data_4;
output 	out_data_buffer_110;
input 	readdata_118;
input 	za_data_11;
input 	readdata_134;
input 	za_data_13;
input 	readdata_164;
input 	readdata_124;
input 	za_data_12;
input 	readdata_57;
input 	za_data_5;
input 	readdata_144;
input 	za_data_14;
input 	readdata_157;
input 	za_data_15;
input 	readdata_104;
input 	za_data_10;
input 	readdata_96;
input 	za_data_9;
input 	readdata_86;
input 	za_data_8;
input 	readdata_77;
input 	za_data_7;
input 	readdata_67;
input 	za_data_6;
input 	readdata_216;
input 	readdata_301;
input 	readdata_291;
input 	readdata_282;
input 	readdata_272;
input 	readdata_262;
input 	readdata_252;
input 	readdata_242;
input 	readdata_234;
input 	readdata_224;
input 	readdata_204;
input 	readdata_194;
input 	readdata_184;
input 	readdata_174;
output 	src_payload25;
input 	read_0;
input 	av_readdata_0;
input 	readdata_010;
input 	av_readdata_9;
output 	src_data_412;
output 	src_data_421;
output 	src_data_431;
output 	src_data_441;
output 	src_data_451;
output 	src_payload26;
input 	av_readdata_1;
input 	readdata_119;
input 	av_readdata_2;
input 	av_readdata_3;
input 	av_readdata_4;
input 	av_readdata_5;
input 	av_readdata_6;
input 	av_readdata_7;
output 	out_data_buffer_210;
output 	src_payload27;
output 	src_data_33;
output 	src_payload28;
output 	src_payload29;
output 	src_data_34;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
output 	src_payload33;
output 	src_payload34;
input 	readdata_312;
output 	src_payload35;
output 	src_payload36;
output 	src_payload37;
output 	src_payload38;
output 	src_payload39;
output 	src_payload40;
output 	src_data_35;
output 	src_payload41;
output 	src_payload42;
output 	src_payload43;
output 	src_payload44;
output 	src_payload45;
output 	src_payload46;
output 	src_payload47;
output 	src_payload48;
output 	src_payload49;
input 	rvalid;
output 	src_payload50;
input 	woverflow;
output 	src_payload51;
output 	src_payload52;
input 	ac;
input 	av_readdata_8;
output 	out_data_buffer_111;
output 	out_data_buffer_32;
output 	src_payload53;
output 	src_payload54;
output 	src_payload55;
output 	src_payload56;
output 	src_payload57;
output 	src_payload58;
output 	src_payload59;
output 	src_payload60;
output 	out_data_buffer_101;
output 	out_data_buffer_41;
output 	out_data_buffer_51;
output 	out_data_buffer_61;
output 	write2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdram_s1_cmd_width_adapter|address_reg[1]~q ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \crosser_001|clock_xer|out_data_buffer[38]~q ;
wire \crosser_003|clock_xer|out_data_buffer[39]~q ;
wire \crosser_001|clock_xer|out_data_buffer[39]~q ;
wire \crosser_003|clock_xer|out_data_buffer[40]~q ;
wire \crosser_001|clock_xer|out_data_buffer[40]~q ;
wire \crosser_001|clock_xer|out_data_buffer[10]~q ;
wire \cpu_data_master_translator|uav_read~0_combout ;
wire \crosser_001|clock_xer|out_data_buffer[0]~q ;
wire \crosser_001|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_001|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \crosser_001|clock_xer|out_valid~combout ;
wire \crosser_003|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_003|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \crosser_003|clock_xer|out_valid~combout ;
wire \epcs_epcs_control_port_translator|wait_latency_counter[0]~q ;
wire \epcs_epcs_control_port_translator|waitrequest_reset_override~q ;
wire \cmd_mux_010|last_cycle~0_combout ;
wire \crosser_003|clock_xer|out_data_buffer[105]~q ;
wire \crosser_001|clock_xer|out_data_buffer[105]~q ;
wire \cmd_mux_010|src_payload[0]~combout ;
wire \crosser_003|clock_xer|out_data_buffer[46]~q ;
wire \crosser_001|clock_xer|out_data_buffer[46]~q ;
wire \crosser_001|clock_xer|out_data_buffer[7]~q ;
wire \port_led_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \router|Equal6~0_combout ;
wire \router|src_channel[12]~0_combout ;
wire \router|Equal2~1_combout ;
wire \router|src_channel[12]~1_combout ;
wire \router|src_channel[12]~3_combout ;
wire \cpu_instruction_master_translator|read_accepted~q ;
wire \cpu_instruction_master_agent|cp_valid~combout ;
wire \router_001|Equal1~4_combout ;
wire \router|Equal5~0_combout ;
wire \router|src_channel[12]~4_combout ;
wire \cpu_instruction_master_translator|uav_read~combout ;
wire \cmd_mux_012|src_data[46]~combout ;
wire \cmd_mux_012|src_data[60]~combout ;
wire \cmd_mux_012|src_data[47]~combout ;
wire \cmd_mux_012|src_data[49]~combout ;
wire \cmd_mux_012|src_data[48]~combout ;
wire \cmd_mux_012|src_data[51]~combout ;
wire \cmd_mux_012|src_data[50]~combout ;
wire \cmd_mux_012|src_data[53]~combout ;
wire \cmd_mux_012|src_data[52]~combout ;
wire \cmd_mux_012|src_data[55]~combout ;
wire \cmd_mux_012|src_data[54]~combout ;
wire \cmd_mux_012|src_data[57]~combout ;
wire \cmd_mux_012|src_data[56]~combout ;
wire \cmd_mux_012|src_data[59]~combout ;
wire \cmd_mux_012|src_data[58]~combout ;
wire \cmd_mux_012|src_data[38]~combout ;
wire \cmd_mux_012|src_data[39]~combout ;
wire \cmd_mux_012|src_data[40]~combout ;
wire \cmd_mux_012|src_data[41]~combout ;
wire \cmd_mux_012|src_data[42]~combout ;
wire \cmd_mux_012|src_data[43]~combout ;
wire \cmd_mux_012|src_data[44]~combout ;
wire \cmd_mux_012|src_data[45]~combout ;
wire \adc_0_adc_slave_translator|read_latency_shift_reg[0]~q ;
wire \crosser_004|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_005|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_005|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \crosser_004|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \crosser_007|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_007|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ;
wire \port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ;
wire \port_sw_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ;
wire \rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg[0]~q ;
wire \rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg[0]~q ;
wire \timer_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \sdram_s1_agent_rdata_fifo|out_valid~q ;
wire \sdram_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][87]~q ;
wire \sdram_s1_agent|rp_valid~combout ;
wire \sdram_s1_agent_rsp_fifo|mem[0][88]~q ;
wire \sdram_s1_agent|uncompressor|burst_uncompress_address_base[1]~q ;
wire \sdram_s1_agent|uncompressor|burst_uncompress_address_offset[1]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][19]~q ;
wire \sdram_s1_agent|comb~0_combout ;
wire \sdram_s1_rsp_width_adapter|always10~1_combout ;
wire \sdram_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][48]~q ;
wire \adc_0_adc_slave_agent|m0_read~0_combout ;
wire \sdram_s1_cmd_width_adapter|count[0]~q ;
wire \cmd_mux_012|last_cycle~0_combout ;
wire \crosser_001|clock_xer|in_ready~0_combout ;
wire \router|src_channel[12]~5_combout ;
wire \cmd_demux|WideOr0~1_combout ;
wire \timer_0_s1_agent|m0_write~1_combout ;
wire \timer_0_s1_translator|read_latency_shift_reg~0_combout ;
wire \rs232_1_avalon_rs232_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \port_key_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \port_gpio_0_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \sys_id_control_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \sys_id_control_slave_translator|wait_latency_counter[1]~q ;
wire \router|always1~0_combout ;
wire \sys_id_control_slave_translator|wait_latency_counter[0]~q ;
wire \cmd_demux|sink_ready~2_combout ;
wire \crosser_002|clock_xer|take_in_data~0_combout ;
wire \router|Equal13~1_combout ;
wire \crosser|clock_xer|in_data_toggle~q ;
wire \crosser|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \cmd_demux|WideOr0~8_combout ;
wire \crosser_003|clock_xer|out_data_buffer[66]~q ;
wire \crosser_001|clock_xer|out_data_buffer[66]~q ;
wire \epcs_epcs_control_port_agent_rsp_fifo|mem_used[0]~q ;
wire \epcs_epcs_control_port_agent_rsp_fifo|mem[0][105]~q ;
wire \epcs_epcs_control_port_translator|read_latency_shift_reg[0]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|mem_used[0]~q ;
wire \epcs_epcs_control_port_agent|rp_valid~0_combout ;
wire \epcs_epcs_control_port_agent_rsp_fifo|mem[0][84]~q ;
wire \epcs_epcs_control_port_agent_rsp_fifo|mem[0][66]~q ;
wire \crosser_006|clock_xer|in_data_toggle~q ;
wire \crosser_006|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \crosser_005|clock_xer|in_data_toggle~q ;
wire \crosser_005|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \crosser_006|clock_xer|take_in_data~0_combout ;
wire \rsp_demux_010|WideOr0~1_combout ;
wire \epcs_epcs_control_port_agent|uncompressor|sink_ready~0_combout ;
wire \crosser_001|clock_xer|out_data_buffer[64]~q ;
wire \epcs_epcs_control_port_agent|nonposted_write_endofpacket~0_combout ;
wire \epcs_epcs_control_port_translator|uav_waitrequest~0_combout ;
wire \crosser_003|clock_xer|take_in_data~2_combout ;
wire \crosser_001|clock_xer|out_data_buffer[6]~q ;
wire \sys_pll_pll_slave_agent_rsp_fifo|mem_used[0]~q ;
wire \crosser_002|clock_xer|out_data_buffer[105]~q ;
wire \crosser_002|clock_xer|out_data_buffer[64]~q ;
wire \sys_pll_pll_slave_agent_rsp_fifo|mem[0][105]~q ;
wire \sys_pll_pll_slave_translator|read_latency_shift_reg[0]~q ;
wire \sys_pll_pll_slave_agent_rdata_fifo|mem_used[0]~q ;
wire \sys_pll_pll_slave_agent|rp_valid~0_combout ;
wire \crosser_007|clock_xer|in_ready~0_combout ;
wire \sys_pll_pll_slave_agent|uncompressor|sink_ready~0_combout ;
wire \cmd_demux|src12_valid~2_combout ;
wire \cmd_mux_012|src_payload[0]~combout ;
wire \sdram_s1_agent|cp_ready~combout ;
wire \cmd_mux_012|src_data[34]~combout ;
wire \cmd_mux_012|src_data[35]~combout ;
wire \crosser_006|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_006|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ;
wire \cmd_mux_009|saved_grant[1]~q ;
wire \port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg~2_combout ;
wire \cpu_debug_mem_slave_agent_rsp_fifo|mem~1_combout ;
wire \cmd_demux_001|src0_valid~0_combout ;
wire \port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg~1_combout ;
wire \port_gpio_0_avalon_parallel_port_slave_translator|read_latency_shift_reg~1_combout ;
wire \rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg~0_combout ;
wire \timer_0_s1_translator|av_waitrequest_generated~0_combout ;
wire \sdram_s1_cmd_width_adapter|out_endofpacket~0_combout ;
wire \sdram_s1_agent_rsp_fifo|mem[0][57]~q ;
wire \sys_id_control_slave_translator|av_waitrequest_generated~1_combout ;
wire \cmd_demux|sink_ready~4_combout ;
wire \sys_id_control_slave_agent|m0_write~0_combout ;
wire \crosser_003|clock_xer|out_data_buffer[84]~q ;
wire \epcs_epcs_control_port_agent|rp_valid~combout ;
wire \crosser_001|clock_xer|out_data_buffer[5]~q ;
wire \sdram_s1_rsp_width_adapter|data_reg[1]~q ;
wire \sdram_s1_rsp_width_adapter|data_reg[3]~q ;
wire \sdram_s1_rsp_width_adapter|data_reg[4]~q ;
wire \router|Equal5~2_combout ;
wire \sys_pll_pll_slave_agent|rp_valid~combout ;
wire \crosser_004|clock_xer|in_data_toggle~q ;
wire \sdram_s1_rsp_width_adapter|data_reg[11]~q ;
wire \sdram_s1_rsp_width_adapter|data_reg[13]~q ;
wire \sdram_s1_rsp_width_adapter|data_reg[5]~q ;
wire \sdram_s1_rsp_width_adapter|data_reg[15]~q ;
wire \crosser_001|clock_xer|out_data_buffer[4]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[0]~q ;
wire \crosser_004|clock_xer|out_valid~combout ;
wire \crosser_005|clock_xer|out_data_buffer[0]~q ;
wire \crosser_004|clock_xer|out_data_buffer[0]~q ;
wire \timer_0_s1_translator|av_readdata_pre[0]~q ;
wire \crosser_007|clock_xer|out_valid~combout ;
wire \crosser_007|clock_xer|out_data_buffer[0]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[1]~q ;
wire \crosser_005|clock_xer|out_data_buffer[1]~q ;
wire \crosser_004|clock_xer|out_data_buffer[1]~q ;
wire \timer_0_s1_translator|av_readdata_pre[1]~q ;
wire \crosser_007|clock_xer|out_data_buffer[1]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[2]~q ;
wire \crosser_005|clock_xer|out_data_buffer[2]~q ;
wire \timer_0_s1_translator|av_readdata_pre[2]~q ;
wire \crosser_004|clock_xer|out_data_buffer[2]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[3]~q ;
wire \crosser_005|clock_xer|out_data_buffer[3]~q ;
wire \timer_0_s1_translator|av_readdata_pre[3]~q ;
wire \crosser_004|clock_xer|out_data_buffer[3]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[4]~q ;
wire \crosser_005|clock_xer|out_data_buffer[4]~q ;
wire \timer_0_s1_translator|av_readdata_pre[4]~q ;
wire \crosser_004|clock_xer|out_data_buffer[4]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[5]~q ;
wire \rsp_demux_009|src0_valid~0_combout ;
wire \crosser_004|clock_xer|out_data_buffer[5]~q ;
wire \timer_0_s1_translator|av_readdata_pre[5]~q ;
wire \crosser_005|clock_xer|out_data_buffer[5]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[6]~q ;
wire \crosser_004|clock_xer|out_data_buffer[6]~q ;
wire \timer_0_s1_translator|av_readdata_pre[6]~q ;
wire \crosser_005|clock_xer|out_data_buffer[6]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[7]~q ;
wire \crosser_004|clock_xer|out_data_buffer[7]~q ;
wire \timer_0_s1_translator|av_readdata_pre[7]~q ;
wire \crosser_005|clock_xer|out_data_buffer[7]~q ;
wire \cmd_mux_012|src_payload~0_combout ;
wire \cmd_mux_012|src_payload~1_combout ;
wire \cmd_mux_012|src_payload~2_combout ;
wire \cmd_mux_012|src_payload~3_combout ;
wire \cmd_mux_012|src_payload~4_combout ;
wire \cmd_mux_012|src_payload~5_combout ;
wire \cmd_mux_012|src_payload~6_combout ;
wire \cmd_mux_012|src_payload~7_combout ;
wire \cmd_mux_012|src_payload~8_combout ;
wire \cmd_mux_012|src_payload~9_combout ;
wire \cmd_mux_012|src_payload~10_combout ;
wire \cmd_mux_012|src_payload~11_combout ;
wire \cmd_mux_012|src_payload~12_combout ;
wire \cmd_mux_012|src_payload~13_combout ;
wire \cmd_mux_012|src_payload~14_combout ;
wire \cmd_mux_012|src_payload~15_combout ;
wire \jtag_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|mem_used[0]~q ;
wire \jtag_avalon_jtag_slave_agent_rsp_fifo|mem[0][105]~q ;
wire \jtag_avalon_jtag_slave_agent_rsp_fifo|mem_used[0]~q ;
wire \jtag_avalon_jtag_slave_agent|rp_valid~combout ;
wire \crosser_004|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \crosser_005|clock_xer|out_data_buffer[23]~q ;
wire \crosser_005|clock_xer|out_data_buffer[22]~q ;
wire \crosser_004|clock_xer|out_data_buffer[22]~q ;
wire \crosser_005|clock_xer|out_data_buffer[21]~q ;
wire \crosser_004|clock_xer|out_data_buffer[21]~q ;
wire \crosser_005|clock_xer|out_data_buffer[20]~q ;
wire \crosser_004|clock_xer|out_data_buffer[20]~q ;
wire \crosser_005|clock_xer|out_data_buffer[19]~q ;
wire \crosser_004|clock_xer|out_data_buffer[19]~q ;
wire \crosser_005|clock_xer|out_data_buffer[18]~q ;
wire \crosser_004|clock_xer|out_data_buffer[18]~q ;
wire \crosser_005|clock_xer|out_data_buffer[17]~q ;
wire \crosser_004|clock_xer|out_data_buffer[17]~q ;
wire \crosser_005|clock_xer|out_data_buffer[16]~q ;
wire \crosser_004|clock_xer|out_data_buffer[16]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[15]~q ;
wire \crosser_004|clock_xer|out_data_buffer[15]~q ;
wire \crosser_005|clock_xer|out_data_buffer[15]~q ;
wire \timer_0_s1_translator|av_readdata_pre[15]~q ;
wire \crosser_004|clock_xer|out_data_buffer[14]~q ;
wire \timer_0_s1_translator|av_readdata_pre[14]~q ;
wire \crosser_005|clock_xer|out_data_buffer[14]~q ;
wire \timer_0_s1_translator|av_readdata_pre[13]~q ;
wire \crosser_005|clock_xer|out_data_buffer[13]~q ;
wire \crosser_004|clock_xer|out_data_buffer[13]~q ;
wire \crosser_004|clock_xer|out_data_buffer[12]~q ;
wire \timer_0_s1_translator|av_readdata_pre[12]~q ;
wire \crosser_005|clock_xer|out_data_buffer[12]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[11]~q ;
wire \timer_0_s1_translator|av_readdata_pre[11]~q ;
wire \crosser_005|clock_xer|out_data_buffer[11]~q ;
wire \timer_0_s1_translator|av_readdata_pre[10]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[10]~q ;
wire \crosser_005|clock_xer|out_data_buffer[10]~q ;
wire \crosser_004|clock_xer|out_data_buffer[10]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[9]~q ;
wire \crosser_004|clock_xer|out_data_buffer[9]~q ;
wire \crosser_005|clock_xer|out_data_buffer[9]~q ;
wire \timer_0_s1_translator|av_readdata_pre[9]~q ;
wire \adc_0_adc_slave_translator|av_readdata_pre[8]~q ;
wire \crosser_004|clock_xer|out_data_buffer[8]~q ;
wire \timer_0_s1_translator|av_readdata_pre[8]~q ;
wire \crosser_005|clock_xer|out_data_buffer[8]~q ;
wire \crosser_001|clock_xer|out_data_buffer[3]~q ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[0]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[0]~0_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[1]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[1]~1_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[2]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[2]~2_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[3]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[3]~3_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[4]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[4]~4_combout ;
wire \jtag_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ;
wire \crosser|clock_xer|out_data_buffer[105]~q ;
wire \crosser|clock_xer|out_data_buffer[64]~q ;
wire \jtag_avalon_jtag_slave_agent|rp_valid~0_combout ;
wire \crosser_004|clock_xer|in_ready~0_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[11]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[11]~5_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[13]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[13]~6_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[16]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[16]~7_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[12]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[12]~8_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[5]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[5]~9_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[14]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[14]~10_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[15]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[15]~11_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[10]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[10]~12_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[9]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[9]~13_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[8]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[8]~14_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[7]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[7]~15_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[6]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[6]~16_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[21]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[21]~17_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[30]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[30]~18_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[29]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[29]~19_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[28]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[28]~20_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[27]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[27]~21_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[26]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[26]~22_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[25]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[25]~23_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[24]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[24]~24_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[23]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[23]~25_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[22]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[22]~26_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[20]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[20]~27_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[19]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[19]~28_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[18]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[18]~29_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[17]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[17]~30_combout ;
wire \crosser_001|clock_xer|out_data_buffer[2]~q ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[0]~0_combout ;
wire \sys_pll_pll_slave_translator|av_readdata_pre[0]~q ;
wire \sys_pll_pll_slave_agent_rdata_fifo|out_data[0]~0_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[1]~1_combout ;
wire \sys_pll_pll_slave_translator|av_readdata_pre[1]~q ;
wire \sys_pll_pll_slave_agent_rdata_fifo|out_data[1]~1_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[2]~2_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[3]~3_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[4]~4_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[5]~5_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[6]~6_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[7]~7_combout ;
wire \epcs_epcs_control_port_translator|av_readdata_pre[31]~q ;
wire \epcs_epcs_control_port_agent_rdata_fifo|out_data[31]~31_combout ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[22]~8_combout ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[21]~9_combout ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[20]~10_combout ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[19]~11_combout ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[18]~12_combout ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[17]~13_combout ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[16]~14_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[15]~15_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[14]~16_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[13]~17_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[12]~18_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[10]~19_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[9]~20_combout ;
wire \jtag_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[8]~21_combout ;
wire \crosser_001|clock_xer|out_data_buffer[1]~q ;
wire \crosser_003|clock_xer|out_data_buffer[41]~q ;
wire \crosser_001|clock_xer|out_data_buffer[41]~q ;
wire \crosser_003|clock_xer|out_data_buffer[42]~q ;
wire \crosser_001|clock_xer|out_data_buffer[42]~q ;
wire \crosser_003|clock_xer|out_data_buffer[43]~q ;
wire \crosser_001|clock_xer|out_data_buffer[43]~q ;
wire \crosser_003|clock_xer|out_data_buffer[44]~q ;
wire \crosser_001|clock_xer|out_data_buffer[44]~q ;
wire \crosser_003|clock_xer|out_data_buffer[45]~q ;
wire \crosser_001|clock_xer|out_data_buffer[45]~q ;
wire \crosser_001|clock_xer|out_data_buffer[11]~q ;
wire \crosser_001|clock_xer|out_data_buffer[13]~q ;
wire \crosser_001|clock_xer|out_data_buffer[12]~q ;
wire \crosser_001|clock_xer|out_data_buffer[14]~q ;
wire \crosser_001|clock_xer|out_data_buffer[15]~q ;
wire \crosser_001|clock_xer|out_data_buffer[9]~q ;
wire \crosser_001|clock_xer|out_data_buffer[8]~q ;
wire \cmd_mux_010|WideOr1~combout ;
wire \cmd_demux_001|src2_valid~2_combout ;
wire \sdram_s1_agent|cp_ready~2_combout ;
wire \rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg~3_combout ;
wire \sdram_s1_agent|rf_source_data[87]~2_combout ;


niosII_altera_merlin_slave_translator_12 sys_pll_pll_slave_translator(
	.wire_pfdena_reg_ena(wire_pfdena_reg_ena),
	.reset(altera_reset_synchronizer_int_chain_out),
	.rst1(rst1),
	.out_data_buffer_66(out_data_buffer_66),
	.read_latency_shift_reg_0(\sys_pll_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\sys_pll_pll_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\sys_pll_pll_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_119,readdata_010}),
	.clk(clk_clk));

niosII_altera_merlin_slave_translator_2 epcs_epcs_control_port_translator(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst1),
	.wait_latency_counter_0(\epcs_epcs_control_port_translator|wait_latency_counter[0]~q ),
	.waitrequest_reset_override1(\epcs_epcs_control_port_translator|waitrequest_reset_override~q ),
	.mem_used_1(mem_used_11),
	.wait_latency_counter_1(wait_latency_counter_1),
	.last_cycle(\cmd_mux_010|last_cycle~0_combout ),
	.src_valid(src_valid),
	.src_valid1(src_valid1),
	.p1_wr_strobe(p1_wr_strobe),
	.src_data_66(src_data_661),
	.av_begintransfer(av_begintransfer),
	.read_latency_shift_reg_0(\epcs_epcs_control_port_translator|read_latency_shift_reg[0]~q ),
	.uav_waitrequest(\epcs_epcs_control_port_translator|uav_waitrequest~0_combout ),
	.av_readdata_pre_0(\epcs_epcs_control_port_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\epcs_epcs_control_port_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\epcs_epcs_control_port_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\epcs_epcs_control_port_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\epcs_epcs_control_port_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_11(\epcs_epcs_control_port_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_13(\epcs_epcs_control_port_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_16(\epcs_epcs_control_port_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_12(\epcs_epcs_control_port_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_5(\epcs_epcs_control_port_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_14(\epcs_epcs_control_port_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\epcs_epcs_control_port_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_10(\epcs_epcs_control_port_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\epcs_epcs_control_port_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_8(\epcs_epcs_control_port_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_7(\epcs_epcs_control_port_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_6(\epcs_epcs_control_port_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_21(\epcs_epcs_control_port_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_30(\epcs_epcs_control_port_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_29(\epcs_epcs_control_port_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_28(\epcs_epcs_control_port_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_27(\epcs_epcs_control_port_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_26(\epcs_epcs_control_port_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_25(\epcs_epcs_control_port_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_24(\epcs_epcs_control_port_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_23(\epcs_epcs_control_port_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_22(\epcs_epcs_control_port_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_20(\epcs_epcs_control_port_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\epcs_epcs_control_port_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\epcs_epcs_control_port_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\epcs_epcs_control_port_translator|av_readdata_pre[17]~q ),
	.av_readdata({readdata_312,readdata_301,readdata_291,readdata_282,readdata_272,readdata_262,readdata_252,readdata_242,readdata_234,readdata_224,readdata_216,readdata_204,readdata_194,readdata_184,readdata_174,readdata_164,readdata_157,readdata_144,readdata_134,readdata_124,readdata_118,
readdata_104,readdata_96,readdata_86,readdata_77,readdata_67,readdata_57,readdata_47,readdata_38,readdata_215,readdata_117,readdata_09}),
	.av_readdata_pre_31(\epcs_epcs_control_port_translator|av_readdata_pre[31]~q ),
	.WideOr1(\cmd_mux_010|WideOr1~combout ));

niosII_altera_merlin_slave_translator_1 cpu_debug_mem_slave_translator(
	.clk(wire_pll7_clk_0),
	.av_readdata({readdata_311,readdata_30,readdata_29,readdata_281,readdata_271,readdata_261,readdata_251,readdata_241,readdata_233,readdata_223,readdata_212,readdata_203,readdata_193,readdata_183,readdata_173,readdata_162,readdata_151,readdata_141,readdata_131,readdata_121,readdata_111,
readdata_10,readdata_9,readdata_8,readdata_74,readdata_64,readdata_54,readdata_4,readdata_3,readdata_2,readdata_12,readdata_06}),
	.reset(r_sync_rst),
	.hold_waitrequest(hold_waitrequest),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.write(\cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.mem(\cpu_debug_mem_slave_agent_rsp_fifo|mem~1_combout ),
	.WideOr1(WideOr12),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_29(av_readdata_pre_29),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_31(av_readdata_pre_31));

niosII_altera_merlin_slave_translator_11 sys_id_control_slave_translator(
	.clk(wire_pll7_clk_0),
	.W_alu_result_3(W_alu_result_3),
	.av_readdata({gnd,W_alu_result_2,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.reset(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.m0_write(m0_write),
	.Equal9(Equal9),
	.Equal6(\router|Equal6~0_combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.mem_used_1(\sys_id_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\sys_id_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\sys_id_control_slave_translator|wait_latency_counter[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.av_waitrequest_generated(\sys_id_control_slave_translator|av_waitrequest_generated~1_combout ),
	.m0_write1(\sys_id_control_slave_agent|m0_write~0_combout ),
	.av_readdata_pre_30(av_readdata_pre_301));

niosII_altera_merlin_slave_translator_9 rs232_1_avalon_rs232_slave_translator(
	.clk(wire_pll7_clk_0),
	.W_alu_result_3(W_alu_result_3),
	.reset(r_sync_rst),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.hold_waitrequest(hold_waitrequest),
	.Equal9(Equal9),
	.Equal6(\router|Equal6~0_combout ),
	.read_latency_shift_reg_0(\rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\rs232_1_avalon_rs232_slave_agent_rsp_fifo|mem_used[1]~q ),
	.read_latency_shift_reg(read_latency_shift_reg1),
	.read_latency_shift_reg1(\rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg~3_combout ));

niosII_altera_merlin_slave_translator_8 rs232_0_avalon_rs232_slave_translator(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.Equal9(Equal9),
	.read_latency_shift_reg_0(\rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(mem_used_14),
	.read_latency_shift_reg(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg~2_combout ),
	.Equal12(Equal121),
	.read_latency_shift_reg1(\rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg2(read_latency_shift_reg3));

niosII_altera_merlin_slave_translator_4 port_gpio_0_avalon_parallel_port_slave_translator(
	.clk(wire_pll7_clk_0),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.reset(r_sync_rst),
	.Equal6(\router|Equal6~0_combout ),
	.src_channel_12(\router|src_channel[12]~1_combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_used_1(\port_gpio_0_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.read_latency_shift_reg(read_latency_shift_reg2),
	.read_latency_shift_reg1(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg~2_combout ),
	.read_latency_shift_reg2(\port_gpio_0_avalon_parallel_port_slave_translator|read_latency_shift_reg~1_combout ));

niosII_altera_merlin_slave_translator_7 port_sw_avalon_parallel_port_slave_translator(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.hold_waitrequest(hold_waitrequest),
	.read_latency_shift_reg_0(\port_sw_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.write(write));

niosII_altera_merlin_slave_translator_5 port_key_avalon_parallel_port_slave_translator(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.hold_waitrequest(hold_waitrequest),
	.read_latency_shift_reg_0(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg~2_combout ),
	.write(write1));

niosII_altera_merlin_slave_translator_6 port_led_avalon_parallel_port_slave_translator(
	.clk(wire_pll7_clk_0),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.reset(r_sync_rst),
	.Equal9(Equal9),
	.mem_used_1(\port_led_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.Equal5(\router|Equal5~0_combout ),
	.read_latency_shift_reg_0(\port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg1(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg~2_combout ),
	.read_latency_shift_reg2(\port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg~1_combout ));

niosII_altera_merlin_slave_translator_3 jtag_avalon_jtag_slave_translator(
	.av_readdata_pre_22(\jtag_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_21(\jtag_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_20(\jtag_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\jtag_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\jtag_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\jtag_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_16(\jtag_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.rst1(rst1),
	.b_full(b_full),
	.out_data_toggle_flopped(out_data_toggle_flopped1),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,av_readdata_7,av_readdata_6,av_readdata_5,av_readdata_4,av_readdata_3,av_readdata_2,av_readdata_1,av_readdata_0}),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.dreg_0(dreg_01),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_16),
	.out_data_buffer_66(out_data_buffer_661),
	.read_latency_shift_reg_0(\jtag_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg(\jtag_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.b_full1(b_full1),
	.counter_reg_bit_21(counter_reg_bit_21),
	.counter_reg_bit_11(counter_reg_bit_11),
	.counter_reg_bit_51(counter_reg_bit_51),
	.counter_reg_bit_41(counter_reg_bit_41),
	.counter_reg_bit_31(counter_reg_bit_31),
	.counter_reg_bit_01(counter_reg_bit_01),
	.av_readdata_pre_0(\jtag_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\jtag_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\jtag_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\jtag_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\jtag_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\jtag_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\jtag_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\jtag_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_15(\jtag_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_14(\jtag_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_13(\jtag_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_12(\jtag_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_10(\jtag_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\jtag_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_8(\jtag_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.read_0(read_0),
	.clk(clk_clk));

niosII_altera_merlin_slave_translator adc_0_adc_slave_translator(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.mem_used_1(mem_used_1),
	.Equal3(Equal3),
	.read_latency_shift_reg_0(\adc_0_adc_slave_translator|read_latency_shift_reg[0]~q ),
	.always0(always0),
	.waitrequest(waitrequest),
	.read_latency_shift_reg(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg~2_combout ),
	.av_readdata_pre_0(\adc_0_adc_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\adc_0_adc_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\adc_0_adc_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\adc_0_adc_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\adc_0_adc_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\adc_0_adc_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\adc_0_adc_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\adc_0_adc_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_15(\adc_0_adc_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_11(\adc_0_adc_slave_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_10(\adc_0_adc_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\adc_0_adc_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_8(\adc_0_adc_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_01(av_readdata_pre_01),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_155,gnd,gnd,gnd,readdata_115,readdata_103,readdata_94,readdata_84,readdata_75,readdata_65,readdata_55,readdata_45,readdata_36,readdata_210,readdata_113,readdata_07}),
	.write(write2));

niosII_altera_merlin_master_translator_1 cpu_instruction_master_translator(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.hold_waitrequest(hold_waitrequest),
	.saved_grant_1(saved_grant_11),
	.i_read(i_read),
	.read_accepted1(\cpu_instruction_master_translator|read_accepted~q ),
	.Equal1(\router_001|Equal1~4_combout ),
	.uav_read1(\cpu_instruction_master_translator|uav_read~combout ),
	.F_pc_9(F_pc_9),
	.last_cycle(\cmd_mux_012|last_cycle~0_combout ),
	.waitrequest(waitrequest1),
	.mem_used_1(mem_used_15),
	.take_in_data(\crosser_003|clock_xer|take_in_data~2_combout ),
	.out_data_toggle_flopped(\crosser_006|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_006|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.src1_valid(src1_valid),
	.read_accepted2(read_accepted1),
	.src1_valid1(src1_valid1),
	.saved_grant_11(\cmd_mux_009|saved_grant[1]~q ));

niosII_altera_merlin_master_translator cpu_data_master_translator(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.d_read(d_read),
	.read_accepted1(read_accepted),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.hold_waitrequest(hold_waitrequest),
	.d_write(d_write),
	.write_accepted1(write_accepted),
	.WideOr1(WideOr11),
	.WideOr0(\cmd_demux|WideOr0~1_combout ),
	.WideOr01(\cmd_demux|WideOr0~8_combout ),
	.av_waitrequest(cpu_data_master_waitrequest),
	.uav_write(uav_write));

niosII_altera_avalon_sc_fifo_4 jtag_avalon_jtag_slave_agent_rdata_fifo(
	.av_readdata_pre_22(\jtag_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_21(\jtag_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_20(\jtag_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\jtag_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\jtag_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\jtag_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_16(\jtag_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.read_latency_shift_reg_0(\jtag_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\jtag_avalon_jtag_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_105_0(\jtag_avalon_jtag_slave_agent_rsp_fifo|mem[0][105]~q ),
	.mem_used_01(\jtag_avalon_jtag_slave_agent_rsp_fifo|mem_used[0]~q ),
	.rp_valid(\jtag_avalon_jtag_slave_agent|rp_valid~0_combout ),
	.in_ready(\crosser_004|clock_xer|in_ready~0_combout ),
	.av_readdata_pre_0(\jtag_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.out_data_0(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[0]~0_combout ),
	.av_readdata_pre_1(\jtag_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.out_data_1(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[1]~1_combout ),
	.av_readdata_pre_2(\jtag_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.out_data_2(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[2]~2_combout ),
	.av_readdata_pre_3(\jtag_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.out_data_3(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[3]~3_combout ),
	.av_readdata_pre_4(\jtag_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.out_data_4(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[4]~4_combout ),
	.av_readdata_pre_5(\jtag_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.out_data_5(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[5]~5_combout ),
	.av_readdata_pre_6(\jtag_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.out_data_6(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[6]~6_combout ),
	.av_readdata_pre_7(\jtag_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.out_data_7(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[7]~7_combout ),
	.out_data_22(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[22]~8_combout ),
	.out_data_21(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[21]~9_combout ),
	.out_data_20(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[20]~10_combout ),
	.out_data_19(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[19]~11_combout ),
	.out_data_18(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[18]~12_combout ),
	.out_data_17(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[17]~13_combout ),
	.out_data_16(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[16]~14_combout ),
	.av_readdata_pre_15(\jtag_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.out_data_15(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[15]~15_combout ),
	.av_readdata_pre_14(\jtag_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.out_data_14(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[14]~16_combout ),
	.av_readdata_pre_13(\jtag_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.out_data_13(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[13]~17_combout ),
	.av_readdata_pre_12(\jtag_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.out_data_12(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[12]~18_combout ),
	.av_readdata_pre_10(\jtag_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.out_data_10(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[10]~19_combout ),
	.av_readdata_pre_9(\jtag_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.out_data_9(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[9]~20_combout ),
	.av_readdata_pre_8(\jtag_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.out_data_8(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[8]~21_combout ),
	.clk(clk_clk));

niosII_altera_avalon_sc_fifo_5 jtag_avalon_jtag_slave_agent_rsp_fifo(
	.reset(altera_reset_synchronizer_int_chain_out),
	.in_data_toggle(\crosser_004|clock_xer|in_data_toggle~q ),
	.out_data_toggle_flopped(out_data_toggle_flopped1),
	.dreg_0(dreg_01),
	.mem_used_1(mem_used_16),
	.out_data_buffer_66(out_data_buffer_661),
	.read_latency_shift_reg_0(\jtag_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\jtag_avalon_jtag_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_105_0(\jtag_avalon_jtag_slave_agent_rsp_fifo|mem[0][105]~q ),
	.mem_used_01(\jtag_avalon_jtag_slave_agent_rsp_fifo|mem_used[0]~q ),
	.dreg_01(\crosser_004|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.out_data_buffer_65(out_data_buffer_652),
	.read_latency_shift_reg(\jtag_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.out_data_buffer_105(\crosser|clock_xer|out_data_buffer[105]~q ),
	.out_data_buffer_64(\crosser|clock_xer|out_data_buffer[64]~q ),
	.in_ready(\crosser_004|clock_xer|in_ready~0_combout ),
	.clk(clk_clk));

niosII_altera_merlin_slave_agent_3 jtag_avalon_jtag_slave_agent(
	.read_latency_shift_reg_0(\jtag_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\jtag_avalon_jtag_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_105_0(\jtag_avalon_jtag_slave_agent_rsp_fifo|mem[0][105]~q ),
	.mem_used_01(\jtag_avalon_jtag_slave_agent_rsp_fifo|mem_used[0]~q ),
	.rp_valid1(\jtag_avalon_jtag_slave_agent|rp_valid~combout ),
	.rp_valid2(\jtag_avalon_jtag_slave_agent|rp_valid~0_combout ));

niosII_altera_avalon_sc_fifo adc_0_adc_slave_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.mem_used_1(mem_used_1),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.hold_waitrequest(hold_waitrequest),
	.Equal3(Equal3),
	.read_latency_shift_reg_0(\adc_0_adc_slave_translator|read_latency_shift_reg[0]~q ),
	.waitrequest(waitrequest),
	.m0_read(\adc_0_adc_slave_agent|m0_read~0_combout ),
	.read_latency_shift_reg(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg~2_combout ));

niosII_altera_merlin_slave_agent adc_0_adc_slave_agent(
	.mem_used_1(mem_used_1),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.Equal3(Equal3),
	.m0_read1(m0_read),
	.m0_read2(\adc_0_adc_slave_agent|m0_read~0_combout ));

niosII_altera_merlin_master_agent_1 cpu_instruction_master_agent(
	.hold_waitrequest(hold_waitrequest),
	.i_read(i_read),
	.read_accepted(\cpu_instruction_master_translator|read_accepted~q ),
	.cp_valid1(\cpu_instruction_master_agent|cp_valid~combout ));

niosII_altera_merlin_master_agent cpu_data_master_agent(
	.clk(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.hold_waitrequest1(hold_waitrequest),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.cp_valid(cp_valid));

niosII_altera_merlin_slave_translator_13 timer_0_s1_translator(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.cp_valid(cp_valid),
	.m0_write(m0_write),
	.Equal4(Equal4),
	.read_latency_shift_reg_0(\timer_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(mem_used_13),
	.m0_write1(\timer_0_s1_agent|m0_write~1_combout ),
	.wait_latency_counter_0(wait_latency_counter_0),
	.wait_latency_counter_1(wait_latency_counter_11),
	.read_latency_shift_reg(\timer_0_s1_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg1(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg~2_combout ),
	.av_waitrequest_generated(\timer_0_s1_translator|av_waitrequest_generated~0_combout ),
	.av_readdata_pre_0(\timer_0_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\timer_0_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\timer_0_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\timer_0_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\timer_0_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\timer_0_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\timer_0_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\timer_0_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_15(\timer_0_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_14(\timer_0_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_13(\timer_0_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_12(\timer_0_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_11(\timer_0_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_10(\timer_0_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\timer_0_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_8(\timer_0_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_156,readdata_143,readdata_133,readdata_123,readdata_116,readdata_102,readdata_95,readdata_85,readdata_76,readdata_66,readdata_56,readdata_46,readdata_37,readdata_214,readdata_114,readdata_08}));

niosII_altera_avalon_sc_fifo_6 port_gpio_0_avalon_parallel_port_slave_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.hold_waitrequest(hold_waitrequest),
	.Equal6(\router|Equal6~0_combout ),
	.src_channel_12(\router|src_channel[12]~1_combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_used_1(\port_gpio_0_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.read_latency_shift_reg(\port_gpio_0_avalon_parallel_port_slave_translator|read_latency_shift_reg~1_combout ));

niosII_altera_avalon_sc_fifo_9 port_sw_avalon_parallel_port_slave_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.reset(r_sync_rst),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.hold_waitrequest(hold_waitrequest),
	.cp_valid(cp_valid),
	.src_channel_12(\router|src_channel[12]~1_combout ),
	.read_latency_shift_reg_0(\port_sw_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.write(write),
	.write1(write2));

niosII_altera_avalon_sc_fifo_7 port_key_avalon_parallel_port_slave_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.reset(r_sync_rst),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.hold_waitrequest(hold_waitrequest),
	.cp_valid(cp_valid),
	.src_channel_12(\router|src_channel[12]~1_combout ),
	.read_latency_shift_reg_0(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\port_key_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.write(write1));

niosII_altera_avalon_sc_fifo_8 port_led_avalon_parallel_port_slave_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.hold_waitrequest(hold_waitrequest),
	.Equal9(Equal9),
	.mem_used_1(\port_led_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.Equal5(\router|Equal5~0_combout ),
	.read_latency_shift_reg_0(\port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg(\port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg~1_combout ));

niosII_niosII_mm_interconnect_0_router_001 router_001(
	.F_pc_24(F_pc_24),
	.F_pc_23(F_pc_23),
	.F_pc_22(F_pc_22),
	.F_pc_21(F_pc_21),
	.F_pc_20(F_pc_20),
	.F_pc_19(F_pc_19),
	.F_pc_18(F_pc_18),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.F_pc_10(F_pc_10),
	.Equal1(\router_001|Equal1~4_combout ));

niosII_niosII_mm_interconnect_0_router router(
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_3(W_alu_result_3),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.Equal3(Equal3),
	.Equal9(Equal9),
	.Equal6(\router|Equal6~0_combout ),
	.src_channel_12(\router|src_channel[12]~0_combout ),
	.Equal2(\router|Equal2~1_combout ),
	.src_channel_121(\router|src_channel[12]~1_combout ),
	.src_channel_122(\router|src_channel[12]~3_combout ),
	.Equal1(Equal1),
	.Equal4(Equal4),
	.Equal5(\router|Equal5~0_combout ),
	.src_channel_123(\router|src_channel[12]~4_combout ),
	.src_channel_124(\router|src_channel[12]~5_combout ),
	.Equal12(Equal12),
	.always1(\router|always1~0_combout ),
	.Equal13(\router|Equal13~1_combout ),
	.Equal121(Equal121),
	.Equal51(\router|Equal5~2_combout ));

niosII_altera_avalon_sc_fifo_17 timer_0_s1_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.hold_waitrequest(hold_waitrequest),
	.Equal4(Equal4),
	.read_latency_shift_reg_0(\timer_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(mem_used_13),
	.wait_latency_counter_1(wait_latency_counter_11),
	.av_waitrequest_generated(\timer_0_s1_translator|av_waitrequest_generated~0_combout ),
	.period_l_wr_strobe(period_l_wr_strobe));

niosII_altera_merlin_slave_agent_13 timer_0_s1_agent(
	.hold_waitrequest(hold_waitrequest),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.m0_write(m0_write),
	.Equal4(Equal4),
	.mem_used_1(mem_used_13),
	.m0_write1(\timer_0_s1_agent|m0_write~1_combout ));

niosII_altera_avalon_sc_fifo_12 sdram_s1_agent_rdata_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.out_valid1(\sdram_s1_agent_rdata_fifo|out_valid~q ),
	.mem_used_0(\sdram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_87_0(\sdram_s1_agent_rsp_fifo|mem[0][87]~q ),
	.out_payload_0(out_payload_0),
	.out_payload_1(out_payload_1),
	.out_payload_2(out_payload_2),
	.out_payload_3(out_payload_3),
	.out_payload_4(out_payload_4),
	.out_payload_11(out_payload_11),
	.out_payload_13(out_payload_13),
	.out_payload_12(out_payload_12),
	.out_payload_5(out_payload_5),
	.out_payload_14(out_payload_14),
	.out_payload_15(out_payload_15),
	.out_payload_10(out_payload_10),
	.out_payload_9(out_payload_9),
	.out_payload_8(out_payload_8),
	.out_payload_7(out_payload_7),
	.out_payload_6(out_payload_6),
	.za_valid(za_valid),
	.za_data_0(za_data_0),
	.za_data_1(za_data_1),
	.za_data_2(za_data_2),
	.za_data_3(za_data_3),
	.za_data_4(za_data_4),
	.za_data_11(za_data_11),
	.za_data_13(za_data_13),
	.za_data_12(za_data_12),
	.za_data_5(za_data_5),
	.za_data_14(za_data_14),
	.za_data_15(za_data_15),
	.za_data_10(za_data_10),
	.za_data_9(za_data_9),
	.za_data_8(za_data_8),
	.za_data_7(za_data_7),
	.za_data_6(za_data_6));

niosII_altera_avalon_sc_fifo_13 sdram_s1_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.address_reg_1(\sdram_s1_cmd_width_adapter|address_reg[1]~q ),
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_01),
	.use_reg(use_reg),
	.saved_grant_1(saved_grant_11),
	.WideOr1(WideOr1),
	.mem_used_7(mem_used_7),
	.src_data_66(src_data_66),
	.out_valid(\sdram_s1_agent_rdata_fifo|out_valid~q ),
	.mem_used_0(\sdram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_87_0(\sdram_s1_agent_rsp_fifo|mem[0][87]~q ),
	.mem_88_0(\sdram_s1_agent_rsp_fifo|mem[0][88]~q ),
	.mem_54_0(mem_54_0),
	.mem_19_0(\sdram_s1_agent_rsp_fifo|mem[0][19]~q ),
	.comb(\sdram_s1_agent|comb~0_combout ),
	.mem_66_0(\sdram_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_48_0(\sdram_s1_agent_rsp_fifo|mem[0][48]~q ),
	.out_endofpacket(\sdram_s1_cmd_width_adapter|out_endofpacket~0_combout ),
	.mem_57_0(\sdram_s1_agent_rsp_fifo|mem[0][57]~q ),
	.cp_ready(\sdram_s1_agent|cp_ready~2_combout ),
	.rf_source_data_87(\sdram_s1_agent|rf_source_data[87]~2_combout ));

niosII_altera_merlin_slave_agent_10 sdram_s1_agent(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.byteen_reg_0(byteen_reg_0),
	.byteen_reg_1(byteen_reg_1),
	.r_sync_rst(r_sync_rst),
	.entries_1(entries_1),
	.entries_0(entries_0),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.d_byteenable_0(d_byteenable_0),
	.saved_grant_0(saved_grant_01),
	.d_byteenable_1(d_byteenable_1),
	.use_reg(use_reg),
	.saved_grant_1(saved_grant_11),
	.WideOr0(WideOr0),
	.Equal0(Equal0),
	.Equal1(Equal1),
	.WideOr1(WideOr1),
	.m0_write1(m0_write1),
	.mem_used_7(mem_used_7),
	.src_data_66(src_data_66),
	.src_valid(src_valid2),
	.src12_valid(src12_valid),
	.m0_write2(m0_write2),
	.out_valid(\sdram_s1_agent_rdata_fifo|out_valid~q ),
	.mem_used_0(\sdram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_87_0(\sdram_s1_agent_rsp_fifo|mem[0][87]~q ),
	.rp_valid1(\sdram_s1_agent|rp_valid~combout ),
	.mem_54_0(mem_54_0),
	.burst_uncompress_address_base_1(\sdram_s1_agent|uncompressor|burst_uncompress_address_base[1]~q ),
	.burst_uncompress_address_offset_1(\sdram_s1_agent|uncompressor|burst_uncompress_address_offset[1]~q ),
	.mem_19_0(\sdram_s1_agent_rsp_fifo|mem[0][19]~q ),
	.comb(\sdram_s1_agent|comb~0_combout ),
	.cp_ready1(\sdram_s1_agent|cp_ready~combout ),
	.mem_57_0(\sdram_s1_agent_rsp_fifo|mem[0][57]~q ),
	.source_addr_1(source_addr_1),
	.cp_ready2(\sdram_s1_agent|cp_ready~2_combout ),
	.rf_source_data_87(\sdram_s1_agent|rf_source_data[87]~2_combout ));

niosII_altera_avalon_sc_fifo_15 sys_pll_pll_slave_agent_rdata_fifo(
	.reset(altera_reset_synchronizer_int_chain_out),
	.mem_used_0(\sys_pll_pll_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_105_0(\sys_pll_pll_slave_agent_rsp_fifo|mem[0][105]~q ),
	.read_latency_shift_reg_0(\sys_pll_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_01(\sys_pll_pll_slave_agent_rdata_fifo|mem_used[0]~q ),
	.rp_valid(\sys_pll_pll_slave_agent|rp_valid~0_combout ),
	.in_ready(\crosser_007|clock_xer|in_ready~0_combout ),
	.av_readdata_pre_0(\sys_pll_pll_slave_translator|av_readdata_pre[0]~q ),
	.out_data_0(\sys_pll_pll_slave_agent_rdata_fifo|out_data[0]~0_combout ),
	.av_readdata_pre_1(\sys_pll_pll_slave_translator|av_readdata_pre[1]~q ),
	.out_data_1(\sys_pll_pll_slave_agent_rdata_fifo|out_data[1]~1_combout ),
	.clk(clk_clk));

niosII_altera_avalon_sc_fifo_16 sys_pll_pll_slave_agent_rsp_fifo(
	.out_data_toggle_flopped(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.mem_used_1(mem_used_12),
	.wire_pfdena_reg_ena(wire_pfdena_reg_ena),
	.out_data_buffer_65(out_data_buffer_651),
	.reset(altera_reset_synchronizer_int_chain_out),
	.rst1(rst1),
	.mem_used_0(\sys_pll_pll_slave_agent_rsp_fifo|mem_used[0]~q ),
	.out_data_buffer_66(out_data_buffer_66),
	.out_data_buffer_105(\crosser_002|clock_xer|out_data_buffer[105]~q ),
	.out_data_buffer_64(\crosser_002|clock_xer|out_data_buffer[64]~q ),
	.mem_105_0(\sys_pll_pll_slave_agent_rsp_fifo|mem[0][105]~q ),
	.sink_ready(\sys_pll_pll_slave_agent|uncompressor|sink_ready~0_combout ),
	.clk(clk_clk));

niosII_altera_merlin_slave_agent_12 sys_pll_pll_slave_agent(
	.mem_used_0(\sys_pll_pll_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_105_0(\sys_pll_pll_slave_agent_rsp_fifo|mem[0][105]~q ),
	.read_latency_shift_reg_0(\sys_pll_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_01(\sys_pll_pll_slave_agent_rdata_fifo|mem_used[0]~q ),
	.rp_valid1(\sys_pll_pll_slave_agent|rp_valid~0_combout ),
	.in_ready(\crosser_007|clock_xer|in_ready~0_combout ),
	.rf_sink_ready(\sys_pll_pll_slave_agent|uncompressor|sink_ready~0_combout ),
	.rp_valid2(\sys_pll_pll_slave_agent|rp_valid~combout ));

niosII_altera_avalon_sc_fifo_2 epcs_epcs_control_port_agent_rdata_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst1),
	.mem_used_0(\epcs_epcs_control_port_agent_rsp_fifo|mem_used[0]~q ),
	.mem_105_0(\epcs_epcs_control_port_agent_rsp_fifo|mem[0][105]~q ),
	.read_latency_shift_reg_0(\epcs_epcs_control_port_translator|read_latency_shift_reg[0]~q ),
	.mem_used_01(\epcs_epcs_control_port_agent_rdata_fifo|mem_used[0]~q ),
	.rp_valid(\epcs_epcs_control_port_agent|rp_valid~0_combout ),
	.WideOr0(\rsp_demux_010|WideOr0~1_combout ),
	.av_readdata_pre_0(\epcs_epcs_control_port_translator|av_readdata_pre[0]~q ),
	.out_data_0(\epcs_epcs_control_port_agent_rdata_fifo|out_data[0]~0_combout ),
	.av_readdata_pre_1(\epcs_epcs_control_port_translator|av_readdata_pre[1]~q ),
	.out_data_1(\epcs_epcs_control_port_agent_rdata_fifo|out_data[1]~1_combout ),
	.av_readdata_pre_2(\epcs_epcs_control_port_translator|av_readdata_pre[2]~q ),
	.out_data_2(\epcs_epcs_control_port_agent_rdata_fifo|out_data[2]~2_combout ),
	.av_readdata_pre_3(\epcs_epcs_control_port_translator|av_readdata_pre[3]~q ),
	.out_data_3(\epcs_epcs_control_port_agent_rdata_fifo|out_data[3]~3_combout ),
	.av_readdata_pre_4(\epcs_epcs_control_port_translator|av_readdata_pre[4]~q ),
	.out_data_4(\epcs_epcs_control_port_agent_rdata_fifo|out_data[4]~4_combout ),
	.av_readdata_pre_11(\epcs_epcs_control_port_translator|av_readdata_pre[11]~q ),
	.out_data_11(\epcs_epcs_control_port_agent_rdata_fifo|out_data[11]~5_combout ),
	.av_readdata_pre_13(\epcs_epcs_control_port_translator|av_readdata_pre[13]~q ),
	.out_data_13(\epcs_epcs_control_port_agent_rdata_fifo|out_data[13]~6_combout ),
	.av_readdata_pre_16(\epcs_epcs_control_port_translator|av_readdata_pre[16]~q ),
	.out_data_16(\epcs_epcs_control_port_agent_rdata_fifo|out_data[16]~7_combout ),
	.av_readdata_pre_12(\epcs_epcs_control_port_translator|av_readdata_pre[12]~q ),
	.out_data_12(\epcs_epcs_control_port_agent_rdata_fifo|out_data[12]~8_combout ),
	.av_readdata_pre_5(\epcs_epcs_control_port_translator|av_readdata_pre[5]~q ),
	.out_data_5(\epcs_epcs_control_port_agent_rdata_fifo|out_data[5]~9_combout ),
	.av_readdata_pre_14(\epcs_epcs_control_port_translator|av_readdata_pre[14]~q ),
	.out_data_14(\epcs_epcs_control_port_agent_rdata_fifo|out_data[14]~10_combout ),
	.av_readdata_pre_15(\epcs_epcs_control_port_translator|av_readdata_pre[15]~q ),
	.out_data_15(\epcs_epcs_control_port_agent_rdata_fifo|out_data[15]~11_combout ),
	.av_readdata_pre_10(\epcs_epcs_control_port_translator|av_readdata_pre[10]~q ),
	.out_data_10(\epcs_epcs_control_port_agent_rdata_fifo|out_data[10]~12_combout ),
	.av_readdata_pre_9(\epcs_epcs_control_port_translator|av_readdata_pre[9]~q ),
	.out_data_9(\epcs_epcs_control_port_agent_rdata_fifo|out_data[9]~13_combout ),
	.av_readdata_pre_8(\epcs_epcs_control_port_translator|av_readdata_pre[8]~q ),
	.out_data_8(\epcs_epcs_control_port_agent_rdata_fifo|out_data[8]~14_combout ),
	.av_readdata_pre_7(\epcs_epcs_control_port_translator|av_readdata_pre[7]~q ),
	.out_data_7(\epcs_epcs_control_port_agent_rdata_fifo|out_data[7]~15_combout ),
	.av_readdata_pre_6(\epcs_epcs_control_port_translator|av_readdata_pre[6]~q ),
	.out_data_6(\epcs_epcs_control_port_agent_rdata_fifo|out_data[6]~16_combout ),
	.av_readdata_pre_21(\epcs_epcs_control_port_translator|av_readdata_pre[21]~q ),
	.out_data_21(\epcs_epcs_control_port_agent_rdata_fifo|out_data[21]~17_combout ),
	.av_readdata_pre_30(\epcs_epcs_control_port_translator|av_readdata_pre[30]~q ),
	.out_data_30(\epcs_epcs_control_port_agent_rdata_fifo|out_data[30]~18_combout ),
	.av_readdata_pre_29(\epcs_epcs_control_port_translator|av_readdata_pre[29]~q ),
	.out_data_29(\epcs_epcs_control_port_agent_rdata_fifo|out_data[29]~19_combout ),
	.av_readdata_pre_28(\epcs_epcs_control_port_translator|av_readdata_pre[28]~q ),
	.out_data_28(\epcs_epcs_control_port_agent_rdata_fifo|out_data[28]~20_combout ),
	.av_readdata_pre_27(\epcs_epcs_control_port_translator|av_readdata_pre[27]~q ),
	.out_data_27(\epcs_epcs_control_port_agent_rdata_fifo|out_data[27]~21_combout ),
	.av_readdata_pre_26(\epcs_epcs_control_port_translator|av_readdata_pre[26]~q ),
	.out_data_26(\epcs_epcs_control_port_agent_rdata_fifo|out_data[26]~22_combout ),
	.av_readdata_pre_25(\epcs_epcs_control_port_translator|av_readdata_pre[25]~q ),
	.out_data_25(\epcs_epcs_control_port_agent_rdata_fifo|out_data[25]~23_combout ),
	.av_readdata_pre_24(\epcs_epcs_control_port_translator|av_readdata_pre[24]~q ),
	.out_data_24(\epcs_epcs_control_port_agent_rdata_fifo|out_data[24]~24_combout ),
	.av_readdata_pre_23(\epcs_epcs_control_port_translator|av_readdata_pre[23]~q ),
	.out_data_23(\epcs_epcs_control_port_agent_rdata_fifo|out_data[23]~25_combout ),
	.av_readdata_pre_22(\epcs_epcs_control_port_translator|av_readdata_pre[22]~q ),
	.out_data_22(\epcs_epcs_control_port_agent_rdata_fifo|out_data[22]~26_combout ),
	.av_readdata_pre_20(\epcs_epcs_control_port_translator|av_readdata_pre[20]~q ),
	.out_data_20(\epcs_epcs_control_port_agent_rdata_fifo|out_data[20]~27_combout ),
	.av_readdata_pre_19(\epcs_epcs_control_port_translator|av_readdata_pre[19]~q ),
	.out_data_19(\epcs_epcs_control_port_agent_rdata_fifo|out_data[19]~28_combout ),
	.av_readdata_pre_18(\epcs_epcs_control_port_translator|av_readdata_pre[18]~q ),
	.out_data_18(\epcs_epcs_control_port_agent_rdata_fifo|out_data[18]~29_combout ),
	.av_readdata_pre_17(\epcs_epcs_control_port_translator|av_readdata_pre[17]~q ),
	.out_data_17(\epcs_epcs_control_port_agent_rdata_fifo|out_data[17]~30_combout ),
	.av_readdata_pre_31(\epcs_epcs_control_port_translator|av_readdata_pre[31]~q ),
	.out_data_31(\epcs_epcs_control_port_agent_rdata_fifo|out_data[31]~31_combout ));

niosII_altera_avalon_sc_fifo_3 epcs_epcs_control_port_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst1),
	.saved_grant_1(saved_grant_1),
	.mem_used_1(mem_used_11),
	.last_cycle(\cmd_mux_010|last_cycle~0_combout ),
	.src_data_66(src_data_661),
	.mem_used_0(\epcs_epcs_control_port_agent_rsp_fifo|mem_used[0]~q ),
	.mem_105_0(\epcs_epcs_control_port_agent_rsp_fifo|mem[0][105]~q ),
	.rp_valid(\epcs_epcs_control_port_agent|rp_valid~0_combout ),
	.mem_84_0(\epcs_epcs_control_port_agent_rsp_fifo|mem[0][84]~q ),
	.mem_66_0(\epcs_epcs_control_port_agent_rsp_fifo|mem[0][66]~q ),
	.WideOr0(\rsp_demux_010|WideOr0~1_combout ),
	.sink_ready(\epcs_epcs_control_port_agent|uncompressor|sink_ready~0_combout ),
	.nonposted_write_endofpacket(\epcs_epcs_control_port_agent|nonposted_write_endofpacket~0_combout ),
	.uav_waitrequest(\epcs_epcs_control_port_translator|uav_waitrequest~0_combout ),
	.out_data_buffer_84(\crosser_003|clock_xer|out_data_buffer[84]~q ),
	.WideOr1(\cmd_mux_010|WideOr1~combout ));

niosII_altera_merlin_slave_agent_2 epcs_epcs_control_port_agent(
	.src_payload_0(\cmd_mux_010|src_payload[0]~combout ),
	.p1_wr_strobe(p1_wr_strobe),
	.mem_used_0(\epcs_epcs_control_port_agent_rsp_fifo|mem_used[0]~q ),
	.mem_105_0(\epcs_epcs_control_port_agent_rsp_fifo|mem[0][105]~q ),
	.read_latency_shift_reg_0(\epcs_epcs_control_port_translator|read_latency_shift_reg[0]~q ),
	.mem_used_01(\epcs_epcs_control_port_agent_rdata_fifo|mem_used[0]~q ),
	.rp_valid1(\epcs_epcs_control_port_agent|rp_valid~0_combout ),
	.WideOr0(\rsp_demux_010|WideOr0~1_combout ),
	.rf_sink_ready(\epcs_epcs_control_port_agent|uncompressor|sink_ready~0_combout ),
	.out_data_buffer_64(\crosser_001|clock_xer|out_data_buffer[64]~q ),
	.nonposted_write_endofpacket(\epcs_epcs_control_port_agent|nonposted_write_endofpacket~0_combout ),
	.rp_valid2(\epcs_epcs_control_port_agent|rp_valid~combout ),
	.WideOr1(\cmd_mux_010|WideOr1~combout ));

niosII_altera_avalon_sc_fifo_1 cpu_debug_mem_slave_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.uav_read1(\cpu_instruction_master_translator|uav_read~combout ),
	.mem_84_0(mem_84_0),
	.mem_66_0(mem_66_0),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.saved_grant_0(saved_grant_02),
	.waitrequest(waitrequest1),
	.mem_used_1(mem_used_15),
	.write(\cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(\cmd_mux_009|saved_grant[1]~q ),
	.mem(\cpu_debug_mem_slave_agent_rsp_fifo|mem~1_combout ),
	.WideOr1(WideOr12),
	.rf_source_valid(rf_source_valid));

niosII_altera_merlin_slave_agent_1 cpu_debug_mem_slave_agent(
	.mem(\cpu_debug_mem_slave_agent_rsp_fifo|mem~1_combout ),
	.WideOr1(WideOr12),
	.rf_source_valid(rf_source_valid));

niosII_altera_avalon_sc_fifo_14 sys_id_control_slave_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.mem_used_1(\sys_id_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.sink_ready1(\cmd_demux|sink_ready~4_combout ));

niosII_altera_merlin_slave_agent_11 sys_id_control_slave_agent(
	.mem_used_1(\sys_id_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.always1(\router|always1~0_combout ),
	.m0_write(\sys_id_control_slave_agent|m0_write~0_combout ));

niosII_altera_avalon_sc_fifo_11 rs232_1_avalon_rs232_slave_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.W_alu_result_3(W_alu_result_3),
	.reset(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.hold_waitrequest(hold_waitrequest),
	.Equal9(Equal9),
	.Equal6(\router|Equal6~0_combout ),
	.read_latency_shift_reg_0(\rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\rs232_1_avalon_rs232_slave_agent_rsp_fifo|mem_used[1]~q ),
	.read_latency_shift_reg(\rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg~3_combout ));

niosII_altera_avalon_sc_fifo_10 rs232_0_avalon_rs232_slave_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg[0]~q ),
	.Equal12(Equal12),
	.mem_used_1(mem_used_14),
	.read_latency_shift_reg(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg~2_combout ),
	.read_latency_shift_reg1(\rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg~0_combout ));

niosII_niosII_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.hold_waitrequest(hold_waitrequest),
	.i_read(i_read),
	.read_accepted(\cpu_instruction_master_translator|read_accepted~q ),
	.Equal1(\router_001|Equal1~4_combout ),
	.uav_read(\cpu_instruction_master_translator|uav_read~combout ),
	.F_pc_9(F_pc_9),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.src2_valid(\cmd_demux_001|src2_valid~2_combout ));

niosII_niosII_mm_interconnect_0_cmd_demux cmd_demux(
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.hold_waitrequest(hold_waitrequest),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.cp_valid(cp_valid),
	.Equal9(Equal9),
	.mem_used_1(\port_led_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_0(saved_grant_01),
	.src_channel_12(\router|src_channel[12]~0_combout ),
	.Equal2(\router|Equal2~1_combout ),
	.src_channel_121(\router|src_channel[12]~1_combout ),
	.src_channel_122(\router|src_channel[12]~3_combout ),
	.Equal1(Equal1),
	.src_channel_123(\router|src_channel[12]~4_combout ),
	.src12_valid(src12_valid),
	.waitrequest(waitrequest),
	.m0_read(\adc_0_adc_slave_agent|m0_read~0_combout ),
	.last_cycle(\cmd_mux_012|last_cycle~0_combout ),
	.in_ready(\crosser_001|clock_xer|in_ready~0_combout ),
	.src_channel_124(\router|src_channel[12]~5_combout ),
	.WideOr0(\cmd_demux|WideOr0~1_combout ),
	.read_latency_shift_reg(\timer_0_s1_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg1(read_latency_shift_reg1),
	.mem_used_11(\port_key_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.mem_used_12(\port_gpio_0_avalon_parallel_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.write(write),
	.Equal12(Equal12),
	.mem_used_13(mem_used_14),
	.mem_used_14(\sys_id_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\sys_id_control_slave_translator|wait_latency_counter[1]~q ),
	.always1(\router|always1~0_combout ),
	.wait_latency_counter_0(\sys_id_control_slave_translator|wait_latency_counter[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.take_in_data(\crosser_002|clock_xer|take_in_data~0_combout ),
	.saved_grant_01(saved_grant_02),
	.waitrequest1(waitrequest1),
	.mem_used_15(mem_used_15),
	.Equal13(\router|Equal13~1_combout ),
	.in_data_toggle(\crosser|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.WideOr01(\cmd_demux|WideOr0~8_combout ),
	.src12_valid1(\cmd_demux|src12_valid~2_combout ),
	.av_waitrequest_generated(\sys_id_control_slave_translator|av_waitrequest_generated~1_combout ),
	.sink_ready1(\cmd_demux|sink_ready~4_combout ));

niosII_altera_avalon_st_handshake_clock_crosser_5 crosser_005(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.r_sync_rst1(r_sync_rst1),
	.out_data_toggle_flopped(\crosser_005|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_005|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.in_data_toggle(\crosser_005|clock_xer|in_data_toggle~q ),
	.dreg_01(\crosser_005|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.take_in_data(\crosser_006|clock_xer|take_in_data~0_combout ),
	.rp_valid(\epcs_epcs_control_port_agent|rp_valid~combout ),
	.out_valid(out_valid1),
	.out_data_buffer_0(\crosser_005|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_1(\crosser_005|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_2(\crosser_005|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_3(\crosser_005|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_4(\crosser_005|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_5(\crosser_005|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_6(\crosser_005|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_7(\crosser_005|clock_xer|out_data_buffer[7]~q ),
	.out_data_buffer_26(out_data_buffer_261),
	.out_data_buffer_25(out_data_buffer_251),
	.out_data_buffer_24(out_data_buffer_241),
	.out_data_buffer_23(\crosser_005|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_22(\crosser_005|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_21(\crosser_005|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_20(\crosser_005|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_19(\crosser_005|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_18(\crosser_005|clock_xer|out_data_buffer[18]~q ),
	.out_data_buffer_17(\crosser_005|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_16(\crosser_005|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_15(\crosser_005|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_14(\crosser_005|clock_xer|out_data_buffer[14]~q ),
	.out_data_buffer_13(\crosser_005|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_12(\crosser_005|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_11(\crosser_005|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_10(\crosser_005|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_9(\crosser_005|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_8(\crosser_005|clock_xer|out_data_buffer[8]~q ),
	.out_data_0(\epcs_epcs_control_port_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\epcs_epcs_control_port_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\epcs_epcs_control_port_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\epcs_epcs_control_port_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\epcs_epcs_control_port_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_buffer_27(out_data_buffer_271),
	.out_data_buffer_28(out_data_buffer_281),
	.out_data_buffer_29(out_data_buffer_291),
	.out_data_buffer_30(out_data_buffer_301),
	.out_data_buffer_31(out_data_buffer_311),
	.out_data_11(\epcs_epcs_control_port_agent_rdata_fifo|out_data[11]~5_combout ),
	.out_data_13(\epcs_epcs_control_port_agent_rdata_fifo|out_data[13]~6_combout ),
	.out_data_16(\epcs_epcs_control_port_agent_rdata_fifo|out_data[16]~7_combout ),
	.out_data_12(\epcs_epcs_control_port_agent_rdata_fifo|out_data[12]~8_combout ),
	.out_data_5(\epcs_epcs_control_port_agent_rdata_fifo|out_data[5]~9_combout ),
	.out_data_14(\epcs_epcs_control_port_agent_rdata_fifo|out_data[14]~10_combout ),
	.out_data_15(\epcs_epcs_control_port_agent_rdata_fifo|out_data[15]~11_combout ),
	.out_data_10(\epcs_epcs_control_port_agent_rdata_fifo|out_data[10]~12_combout ),
	.out_data_9(\epcs_epcs_control_port_agent_rdata_fifo|out_data[9]~13_combout ),
	.out_data_8(\epcs_epcs_control_port_agent_rdata_fifo|out_data[8]~14_combout ),
	.out_data_7(\epcs_epcs_control_port_agent_rdata_fifo|out_data[7]~15_combout ),
	.out_data_6(\epcs_epcs_control_port_agent_rdata_fifo|out_data[6]~16_combout ),
	.out_data_21(\epcs_epcs_control_port_agent_rdata_fifo|out_data[21]~17_combout ),
	.out_data_30(\epcs_epcs_control_port_agent_rdata_fifo|out_data[30]~18_combout ),
	.out_data_29(\epcs_epcs_control_port_agent_rdata_fifo|out_data[29]~19_combout ),
	.out_data_28(\epcs_epcs_control_port_agent_rdata_fifo|out_data[28]~20_combout ),
	.out_data_27(\epcs_epcs_control_port_agent_rdata_fifo|out_data[27]~21_combout ),
	.out_data_26(\epcs_epcs_control_port_agent_rdata_fifo|out_data[26]~22_combout ),
	.out_data_25(\epcs_epcs_control_port_agent_rdata_fifo|out_data[25]~23_combout ),
	.out_data_24(\epcs_epcs_control_port_agent_rdata_fifo|out_data[24]~24_combout ),
	.out_data_23(\epcs_epcs_control_port_agent_rdata_fifo|out_data[23]~25_combout ),
	.out_data_22(\epcs_epcs_control_port_agent_rdata_fifo|out_data[22]~26_combout ),
	.out_data_20(\epcs_epcs_control_port_agent_rdata_fifo|out_data[20]~27_combout ),
	.out_data_19(\epcs_epcs_control_port_agent_rdata_fifo|out_data[19]~28_combout ),
	.out_data_18(\epcs_epcs_control_port_agent_rdata_fifo|out_data[18]~29_combout ),
	.out_data_17(\epcs_epcs_control_port_agent_rdata_fifo|out_data[17]~30_combout ),
	.out_data_31(\epcs_epcs_control_port_agent_rdata_fifo|out_data[31]~31_combout ));

niosII_altera_avalon_st_handshake_clock_crosser_4 crosser_004(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.out_data_toggle_flopped(\crosser_004|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_004|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.in_data_toggle(\crosser_004|clock_xer|in_data_toggle~q ),
	.out_valid(\crosser_004|clock_xer|out_valid~combout ),
	.out_data_buffer_0(\crosser_004|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_1(\crosser_004|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_2(\crosser_004|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_3(\crosser_004|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_4(\crosser_004|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_5(\crosser_004|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_6(\crosser_004|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_7(\crosser_004|clock_xer|out_data_buffer[7]~q ),
	.rp_valid(\jtag_avalon_jtag_slave_agent|rp_valid~combout ),
	.dreg_01(\crosser_004|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.out_data_buffer_22(\crosser_004|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_21(\crosser_004|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_20(\crosser_004|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_19(\crosser_004|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_18(\crosser_004|clock_xer|out_data_buffer[18]~q ),
	.out_data_buffer_17(\crosser_004|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_16(\crosser_004|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_15(\crosser_004|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_14(\crosser_004|clock_xer|out_data_buffer[14]~q ),
	.out_data_buffer_13(\crosser_004|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_12(\crosser_004|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_10(\crosser_004|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_9(\crosser_004|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_8(\crosser_004|clock_xer|out_data_buffer[8]~q ),
	.in_ready(\crosser_004|clock_xer|in_ready~0_combout ),
	.out_data_0(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_5(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[5]~5_combout ),
	.out_data_6(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[6]~6_combout ),
	.out_data_7(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[7]~7_combout ),
	.out_data_22(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[22]~8_combout ),
	.out_data_21(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[21]~9_combout ),
	.out_data_20(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[20]~10_combout ),
	.out_data_19(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[19]~11_combout ),
	.out_data_18(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[18]~12_combout ),
	.out_data_17(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[17]~13_combout ),
	.out_data_16(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[16]~14_combout ),
	.out_data_15(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[15]~15_combout ),
	.out_data_14(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[14]~16_combout ),
	.out_data_13(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[13]~17_combout ),
	.out_data_12(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[12]~18_combout ),
	.out_data_10(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[10]~19_combout ),
	.out_data_9(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[9]~20_combout ),
	.out_data_8(\jtag_avalon_jtag_slave_agent_rdata_fifo|out_data[8]~21_combout ),
	.clk_clk(clk_clk));

niosII_altera_avalon_st_handshake_clock_crosser_3 crosser_003(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.r_sync_rst1(r_sync_rst1),
	.saved_grant_1(saved_grant_1),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(\crosser_003|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_40(\crosser_003|clock_xer|out_data_buffer[40]~q ),
	.hold_waitrequest(hold_waitrequest),
	.out_data_toggle_flopped(\crosser_003|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_003|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(\crosser_003|clock_xer|out_valid~combout ),
	.last_cycle(\cmd_mux_010|last_cycle~0_combout ),
	.out_data_buffer_105(\crosser_003|clock_xer|out_data_buffer[105]~q ),
	.out_data_buffer_46(\crosser_003|clock_xer|out_data_buffer[46]~q ),
	.i_read(i_read),
	.read_accepted(\cpu_instruction_master_translator|read_accepted~q ),
	.cp_valid(\cpu_instruction_master_agent|cp_valid~combout ),
	.Equal1(\router_001|Equal1~4_combout ),
	.uav_read(\cpu_instruction_master_translator|uav_read~combout ),
	.F_pc_8(F_pc_8),
	.F_pc_9(F_pc_9),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_7(F_pc_7),
	.out_data_buffer_66(\crosser_003|clock_xer|out_data_buffer[66]~q ),
	.take_in_data(\crosser_003|clock_xer|take_in_data~2_combout ),
	.out_data_buffer_84(\crosser_003|clock_xer|out_data_buffer[84]~q ),
	.out_data_buffer_41(\crosser_003|clock_xer|out_data_buffer[41]~q ),
	.out_data_buffer_42(\crosser_003|clock_xer|out_data_buffer[42]~q ),
	.out_data_buffer_43(\crosser_003|clock_xer|out_data_buffer[43]~q ),
	.out_data_buffer_44(\crosser_003|clock_xer|out_data_buffer[44]~q ),
	.out_data_buffer_45(\crosser_003|clock_xer|out_data_buffer[45]~q ));

niosII_altera_avalon_st_handshake_clock_crosser_2 crosser_002(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.r_sync_rst(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.d_writedata_0(d_writedata_0),
	.d_writedata_1(d_writedata_1),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_toggle_flopped(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.mem_used_1(mem_used_12),
	.out_data_buffer_65(out_data_buffer_651),
	.out_data_buffer_38(out_data_buffer_381),
	.out_data_buffer_39(out_data_buffer_39),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_channel_12(\router|src_channel[12]~1_combout ),
	.Equal5(\router|Equal5~0_combout ),
	.take_in_data(\crosser_002|clock_xer|take_in_data~0_combout ),
	.rst1(rst1),
	.out_data_buffer_66(out_data_buffer_66),
	.out_data_buffer_105(\crosser_002|clock_xer|out_data_buffer[105]~q ),
	.out_data_buffer_64(\crosser_002|clock_xer|out_data_buffer[64]~q ),
	.uav_write(uav_write),
	.Equal51(\router|Equal5~2_combout ),
	.out_data_buffer_1(out_data_buffer_111),
	.clk_clk(clk_clk));

niosII_altera_avalon_st_handshake_clock_crosser_1 crosser_001(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.r_sync_rst(r_sync_rst),
	.r_sync_rst1(r_sync_rst1),
	.saved_grant_0(saved_grant_0),
	.out_data_buffer_38(\crosser_001|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_39(\crosser_001|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_40(\crosser_001|clock_xer|out_data_buffer[40]~q ),
	.out_data_buffer_10(\crosser_001|clock_xer|out_data_buffer[10]~q ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.out_data_buffer_0(\crosser_001|clock_xer|out_data_buffer[0]~q ),
	.out_data_toggle_flopped(\crosser_001|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_001|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(\crosser_001|clock_xer|out_valid~combout ),
	.last_cycle(\cmd_mux_010|last_cycle~0_combout ),
	.out_data_buffer_105(\crosser_001|clock_xer|out_data_buffer[105]~q ),
	.out_data_buffer_46(\crosser_001|clock_xer|out_data_buffer[46]~q ),
	.out_data_buffer_65(out_data_buffer_65),
	.out_data_buffer_7(\crosser_001|clock_xer|out_data_buffer[7]~q ),
	.d_writedata_0(d_writedata_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.Equal1(Equal1),
	.src12_valid(src12_valid),
	.in_ready(\crosser_001|clock_xer|in_ready~0_combout ),
	.out_data_buffer_66(\crosser_001|clock_xer|out_data_buffer[66]~q ),
	.out_data_buffer_64(\crosser_001|clock_xer|out_data_buffer[64]~q ),
	.d_writedata_10(d_writedata_10),
	.out_data_buffer_6(\crosser_001|clock_xer|out_data_buffer[6]~q ),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.uav_write(uav_write),
	.out_data_buffer_5(\crosser_001|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_4(\crosser_001|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_3(\crosser_001|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_2(\crosser_001|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_1(\crosser_001|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_41(\crosser_001|clock_xer|out_data_buffer[41]~q ),
	.out_data_buffer_42(\crosser_001|clock_xer|out_data_buffer[42]~q ),
	.out_data_buffer_43(\crosser_001|clock_xer|out_data_buffer[43]~q ),
	.out_data_buffer_44(\crosser_001|clock_xer|out_data_buffer[44]~q ),
	.out_data_buffer_45(\crosser_001|clock_xer|out_data_buffer[45]~q ),
	.out_data_buffer_11(\crosser_001|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_13(\crosser_001|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_12(\crosser_001|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_14(\crosser_001|clock_xer|out_data_buffer[14]~q ),
	.out_data_buffer_15(\crosser_001|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_9(\crosser_001|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_8(\crosser_001|clock_xer|out_data_buffer[8]~q ));

niosII_altera_avalon_st_handshake_clock_crosser crosser(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.W_alu_result_2(W_alu_result_2),
	.r_sync_rst(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.d_writedata_0(d_writedata_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal13(\router|Equal13~1_combout ),
	.in_data_toggle(\crosser|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.d_writedata_10(d_writedata_10),
	.uav_write(uav_write),
	.out_data_toggle_flopped(out_data_toggle_flopped1),
	.dreg_01(dreg_01),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_16),
	.out_data_buffer_66(out_data_buffer_661),
	.out_data_buffer_38(out_data_buffer_382),
	.out_data_buffer_7(out_data_buffer_71),
	.out_data_buffer_65(out_data_buffer_652),
	.out_data_buffer_105(\crosser|clock_xer|out_data_buffer[105]~q ),
	.out_data_buffer_64(\crosser|clock_xer|out_data_buffer[64]~q ),
	.out_data_buffer_0(out_data_buffer_02),
	.out_data_buffer_1(out_data_buffer_110),
	.out_data_buffer_2(out_data_buffer_210),
	.out_data_buffer_3(out_data_buffer_32),
	.out_data_buffer_10(out_data_buffer_101),
	.out_data_buffer_4(out_data_buffer_41),
	.out_data_buffer_5(out_data_buffer_51),
	.out_data_buffer_6(out_data_buffer_61),
	.clk_clk(clk_clk));

niosII_altera_merlin_width_adapter sdram_s1_cmd_width_adapter(
	.clk(wire_pll7_clk_0),
	.byteen_reg_0(byteen_reg_0),
	.byteen_reg_1(byteen_reg_1),
	.address_reg_1(\sdram_s1_cmd_width_adapter|address_reg[1]~q ),
	.reset(r_sync_rst),
	.d_writedata_0(d_writedata_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.saved_grant_0(saved_grant_01),
	.use_reg1(use_reg),
	.WideOr0(WideOr0),
	.Equal0(Equal0),
	.WideOr1(WideOr1),
	.mem_used_7(mem_used_7),
	.src_data_46(\cmd_mux_012|src_data[46]~combout ),
	.out_data_28(out_data_28),
	.src_data_60(\cmd_mux_012|src_data[60]~combout ),
	.out_data_42(out_data_42),
	.src_data_47(\cmd_mux_012|src_data[47]~combout ),
	.out_data_29(out_data_29),
	.src_data_49(\cmd_mux_012|src_data[49]~combout ),
	.out_data_31(out_data_31),
	.src_data_48(\cmd_mux_012|src_data[48]~combout ),
	.out_data_30(out_data_30),
	.src_data_51(\cmd_mux_012|src_data[51]~combout ),
	.out_data_33(out_data_33),
	.src_data_50(\cmd_mux_012|src_data[50]~combout ),
	.out_data_32(out_data_32),
	.src_data_53(\cmd_mux_012|src_data[53]~combout ),
	.out_data_35(out_data_35),
	.src_data_52(\cmd_mux_012|src_data[52]~combout ),
	.out_data_34(out_data_34),
	.src_data_55(\cmd_mux_012|src_data[55]~combout ),
	.out_data_37(out_data_37),
	.src_data_54(\cmd_mux_012|src_data[54]~combout ),
	.out_data_36(out_data_36),
	.src_data_57(\cmd_mux_012|src_data[57]~combout ),
	.out_data_39(out_data_39),
	.src_data_56(\cmd_mux_012|src_data[56]~combout ),
	.out_data_38(out_data_38),
	.src_data_59(\cmd_mux_012|src_data[59]~combout ),
	.out_data_41(out_data_41),
	.src_data_58(\cmd_mux_012|src_data[58]~combout ),
	.out_data_40(out_data_40),
	.out_data_19(out_data_19),
	.src_data_38(\cmd_mux_012|src_data[38]~combout ),
	.out_data_20(out_data_20),
	.src_data_39(\cmd_mux_012|src_data[39]~combout ),
	.out_data_21(out_data_21),
	.src_data_40(\cmd_mux_012|src_data[40]~combout ),
	.out_data_22(out_data_22),
	.src_data_41(\cmd_mux_012|src_data[41]~combout ),
	.out_data_23(out_data_23),
	.src_data_42(\cmd_mux_012|src_data[42]~combout ),
	.out_data_24(out_data_24),
	.src_data_43(\cmd_mux_012|src_data[43]~combout ),
	.out_data_25(out_data_25),
	.src_data_44(\cmd_mux_012|src_data[44]~combout ),
	.out_data_26(out_data_26),
	.src_data_45(\cmd_mux_012|src_data[45]~combout ),
	.out_data_27(out_data_27),
	.count_0(\sdram_s1_cmd_width_adapter|count[0]~q ),
	.d_writedata_10(d_writedata_10),
	.in_endofpacket(\cmd_mux_012|src_payload[0]~combout ),
	.cp_ready(\sdram_s1_agent|cp_ready~combout ),
	.src_data_34(\cmd_mux_012|src_data[34]~combout ),
	.src_data_35(\cmd_mux_012|src_data[35]~combout ),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.out_endofpacket(\sdram_s1_cmd_width_adapter|out_endofpacket~0_combout ),
	.out_data_0(out_data_0),
	.out_data_1(out_data_1),
	.out_data_2(out_data_2),
	.out_data_3(out_data_3),
	.out_data_4(out_data_4),
	.out_data_5(out_data_5),
	.out_data_6(out_data_6),
	.out_data_7(out_data_7),
	.out_data_8(out_data_8),
	.out_data_9(out_data_9),
	.out_data_10(out_data_10),
	.out_data_11(out_data_11),
	.out_data_12(out_data_12),
	.out_data_13(out_data_13),
	.out_data_14(out_data_14),
	.out_data_15(out_data_15),
	.src_payload(\cmd_mux_012|src_payload~0_combout ),
	.src_payload1(\cmd_mux_012|src_payload~1_combout ),
	.src_payload2(\cmd_mux_012|src_payload~2_combout ),
	.src_payload3(\cmd_mux_012|src_payload~3_combout ),
	.src_payload4(\cmd_mux_012|src_payload~4_combout ),
	.src_payload5(\cmd_mux_012|src_payload~5_combout ),
	.src_payload6(\cmd_mux_012|src_payload~6_combout ),
	.src_payload7(\cmd_mux_012|src_payload~7_combout ),
	.src_payload8(\cmd_mux_012|src_payload~8_combout ),
	.src_payload9(\cmd_mux_012|src_payload~9_combout ),
	.src_payload10(\cmd_mux_012|src_payload~10_combout ),
	.src_payload11(\cmd_mux_012|src_payload~11_combout ),
	.src_payload12(\cmd_mux_012|src_payload~12_combout ),
	.src_payload13(\cmd_mux_012|src_payload~13_combout ),
	.src_payload14(\cmd_mux_012|src_payload~14_combout ),
	.src_payload15(\cmd_mux_012|src_payload~15_combout ));

niosII_altera_merlin_width_adapter_1 sdram_s1_rsp_width_adapter(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.rp_valid(\sdram_s1_agent|rp_valid~combout ),
	.mem_88_0(\sdram_s1_agent_rsp_fifo|mem[0][88]~q ),
	.mem_54_0(mem_54_0),
	.burst_uncompress_address_base_1(\sdram_s1_agent|uncompressor|burst_uncompress_address_base[1]~q ),
	.burst_uncompress_address_offset_1(\sdram_s1_agent|uncompressor|burst_uncompress_address_offset[1]~q ),
	.mem_19_0(\sdram_s1_agent_rsp_fifo|mem[0][19]~q ),
	.comb(\sdram_s1_agent|comb~0_combout ),
	.always10(\sdram_s1_rsp_width_adapter|always10~1_combout ),
	.data_reg_0(data_reg_0),
	.out_payload_0(out_payload_0),
	.source_addr_1(source_addr_1),
	.data_reg_1(\sdram_s1_rsp_width_adapter|data_reg[1]~q ),
	.out_payload_1(out_payload_1),
	.data_reg_2(data_reg_2),
	.out_payload_2(out_payload_2),
	.data_reg_3(\sdram_s1_rsp_width_adapter|data_reg[3]~q ),
	.out_payload_3(out_payload_3),
	.data_reg_4(\sdram_s1_rsp_width_adapter|data_reg[4]~q ),
	.out_payload_4(out_payload_4),
	.data_reg_11(\sdram_s1_rsp_width_adapter|data_reg[11]~q ),
	.out_payload_11(out_payload_11),
	.data_reg_13(\sdram_s1_rsp_width_adapter|data_reg[13]~q ),
	.out_payload_13(out_payload_13),
	.data_reg_12(data_reg_12),
	.out_payload_12(out_payload_12),
	.data_reg_5(\sdram_s1_rsp_width_adapter|data_reg[5]~q ),
	.out_payload_5(out_payload_5),
	.data_reg_14(data_reg_14),
	.out_payload_14(out_payload_14),
	.data_reg_15(\sdram_s1_rsp_width_adapter|data_reg[15]~q ),
	.out_payload_15(out_payload_15),
	.data_reg_10(data_reg_10),
	.out_payload_10(out_payload_10),
	.data_reg_9(data_reg_9),
	.out_payload_9(out_payload_9),
	.data_reg_8(data_reg_8),
	.out_payload_8(out_payload_8),
	.data_reg_7(data_reg_7),
	.out_payload_7(out_payload_7),
	.data_reg_6(data_reg_6),
	.out_payload_6(out_payload_6));

niosII_niosII_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.src1_valid(src1_valid1),
	.source_addr_1(source_addr_1),
	.src_payload(src_payload6));

niosII_niosII_mm_interconnect_0_rsp_mux rsp_mux(
	.readdata_0(readdata_0),
	.readdata_01(readdata_01),
	.readdata_1(readdata_1),
	.readdata_11(readdata_11),
	.readdata_23(readdata_23),
	.readdata_231(readdata_231),
	.readdata_22(readdata_22),
	.readdata_221(readdata_221),
	.readdata_21(readdata_21),
	.readdata_211(readdata_211),
	.readdata_20(readdata_20),
	.readdata_201(readdata_201),
	.readdata_19(readdata_19),
	.readdata_191(readdata_191),
	.readdata_18(readdata_18),
	.readdata_181(readdata_181),
	.readdata_17(readdata_17),
	.readdata_171(readdata_171),
	.readdata_16(readdata_16),
	.readdata_161(readdata_161),
	.read_latency_shift_reg_0(\adc_0_adc_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_84_0(mem_84_0),
	.mem_66_0(mem_66_0),
	.read_latency_shift_reg_01(read_latency_shift_reg_0),
	.out_data_toggle_flopped(\crosser_004|clock_xer|out_data_toggle_flopped~q ),
	.out_data_toggle_flopped1(\crosser_005|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_005|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.dreg_01(\crosser_004|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_data_toggle_flopped2(\crosser_007|clock_xer|out_data_toggle_flopped~q ),
	.dreg_02(\crosser_007|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.read_latency_shift_reg_02(\port_led_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\port_key_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_04(\port_sw_avalon_parallel_port_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_05(read_latency_shift_reg_01),
	.read_latency_shift_reg_06(\rs232_0_avalon_rs232_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_07(\rs232_1_avalon_rs232_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_08(read_latency_shift_reg_02),
	.read_latency_shift_reg_09(\timer_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_54_0(mem_54_0),
	.src0_valid(src0_valid),
	.WideOr11(WideOr11),
	.av_readdata_pre_0(av_readdata_pre_0),
	.out_payload_0(out_payload_0),
	.source_addr_1(source_addr_1),
	.F_iw_0(F_iw_0),
	.av_readdata_pre_1(av_readdata_pre_1),
	.data_reg_1(\sdram_s1_rsp_width_adapter|data_reg[1]~q ),
	.out_payload_1(out_payload_1),
	.src_data_1(src_data_1),
	.av_readdata_pre_2(av_readdata_pre_2),
	.out_payload_2(out_payload_2),
	.F_iw_2(F_iw_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.data_reg_3(\sdram_s1_rsp_width_adapter|data_reg[3]~q ),
	.out_payload_3(out_payload_3),
	.src_data_3(src_data_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.data_reg_4(\sdram_s1_rsp_width_adapter|data_reg[4]~q ),
	.out_payload_4(out_payload_4),
	.src_data_4(src_data_4),
	.av_readdata_pre_11(av_readdata_pre_11),
	.data_reg_11(\sdram_s1_rsp_width_adapter|data_reg[11]~q ),
	.out_payload_11(out_payload_11),
	.src_data_11(src_data_11),
	.av_readdata_pre_13(av_readdata_pre_13),
	.data_reg_13(\sdram_s1_rsp_width_adapter|data_reg[13]~q ),
	.out_payload_13(out_payload_13),
	.src_data_13(src_data_13),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.F_iw_12(F_iw_12),
	.av_readdata_pre_5(av_readdata_pre_5),
	.data_reg_5(\sdram_s1_rsp_width_adapter|data_reg[5]~q ),
	.out_payload_5(out_payload_5),
	.src_data_5(src_data_5),
	.av_readdata_pre_14(av_readdata_pre_14),
	.F_iw_14(F_iw_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.data_reg_15(\sdram_s1_rsp_width_adapter|data_reg[15]~q ),
	.out_payload_15(out_payload_15),
	.src_data_15(src_data_15),
	.av_readdata_pre_10(av_readdata_pre_10),
	.F_iw_10(F_iw_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.F_iw_9(F_iw_9),
	.av_readdata_pre_8(av_readdata_pre_8),
	.F_iw_8(F_iw_8),
	.av_readdata_pre_7(av_readdata_pre_7),
	.out_payload_7(out_payload_7),
	.F_iw_7(F_iw_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.out_payload_6(out_payload_6),
	.F_iw_6(F_iw_6),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.readdata_02(readdata_02),
	.av_readdata_pre_01(\adc_0_adc_slave_translator|av_readdata_pre[0]~q ),
	.readdata_03(readdata_03),
	.readdata_04(readdata_04),
	.readdata_05(readdata_05),
	.out_valid(\crosser_004|clock_xer|out_valid~combout ),
	.out_valid1(out_valid1),
	.out_data_buffer_0(\crosser_005|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_01(\crosser_004|clock_xer|out_data_buffer[0]~q ),
	.av_readdata_pre_02(\timer_0_s1_translator|av_readdata_pre[0]~q ),
	.out_valid2(\crosser_007|clock_xer|out_valid~combout ),
	.out_data_buffer_02(\crosser_007|clock_xer|out_data_buffer[0]~q ),
	.src_data_0(src_data_0),
	.readdata_12(readdata_13),
	.av_readdata_pre_110(\adc_0_adc_slave_translator|av_readdata_pre[1]~q ),
	.readdata_13(readdata_14),
	.readdata_14(readdata_15),
	.readdata_15(readdata_110),
	.out_data_buffer_1(\crosser_005|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_11(\crosser_004|clock_xer|out_data_buffer[1]~q ),
	.av_readdata_pre_111(\timer_0_s1_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_12(\crosser_007|clock_xer|out_data_buffer[1]~q ),
	.src_data_12(src_data_12),
	.src_data_2(src_data_2),
	.readdata_2(readdata_24),
	.av_readdata_pre_24(\adc_0_adc_slave_translator|av_readdata_pre[2]~q ),
	.readdata_24(readdata_25),
	.readdata_25(readdata_26),
	.readdata_26(readdata_27),
	.readdata_27(readdata_28),
	.out_data_buffer_2(\crosser_005|clock_xer|out_data_buffer[2]~q ),
	.av_readdata_pre_25(\timer_0_s1_translator|av_readdata_pre[2]~q ),
	.out_data_buffer_21(\crosser_004|clock_xer|out_data_buffer[2]~q ),
	.src_data_21(src_data_21),
	.readdata_3(readdata_31),
	.av_readdata_pre_31(\adc_0_adc_slave_translator|av_readdata_pre[3]~q ),
	.readdata_31(readdata_32),
	.readdata_32(readdata_33),
	.readdata_33(readdata_34),
	.readdata_34(readdata_35),
	.out_data_buffer_3(\crosser_005|clock_xer|out_data_buffer[3]~q ),
	.av_readdata_pre_32(\timer_0_s1_translator|av_readdata_pre[3]~q ),
	.out_data_buffer_31(\crosser_004|clock_xer|out_data_buffer[3]~q ),
	.src_data_31(src_data_31),
	.readdata_4(readdata_41),
	.av_readdata_pre_41(\adc_0_adc_slave_translator|av_readdata_pre[4]~q ),
	.readdata_41(readdata_42),
	.readdata_42(readdata_43),
	.readdata_43(readdata_44),
	.av_readdata_pre_30(av_readdata_pre_301),
	.out_data_buffer_4(\crosser_005|clock_xer|out_data_buffer[4]~q ),
	.av_readdata_pre_42(\timer_0_s1_translator|av_readdata_pre[4]~q ),
	.out_data_buffer_41(\crosser_004|clock_xer|out_data_buffer[4]~q ),
	.src_data_41(src_data_41),
	.readdata_5(readdata_5),
	.av_readdata_pre_51(\adc_0_adc_slave_translator|av_readdata_pre[5]~q ),
	.src0_valid1(\rsp_demux_009|src0_valid~0_combout ),
	.readdata_51(readdata_51),
	.readdata_52(readdata_52),
	.out_data_buffer_5(\crosser_004|clock_xer|out_data_buffer[5]~q ),
	.readdata_53(readdata_53),
	.av_readdata_pre_52(\timer_0_s1_translator|av_readdata_pre[5]~q ),
	.out_data_buffer_51(\crosser_005|clock_xer|out_data_buffer[5]~q ),
	.src_data_51(src_data_51),
	.readdata_6(readdata_6),
	.av_readdata_pre_61(\adc_0_adc_slave_translator|av_readdata_pre[6]~q ),
	.readdata_61(readdata_61),
	.readdata_62(readdata_62),
	.out_data_buffer_6(\crosser_004|clock_xer|out_data_buffer[6]~q ),
	.readdata_63(readdata_63),
	.av_readdata_pre_62(\timer_0_s1_translator|av_readdata_pre[6]~q ),
	.out_data_buffer_61(\crosser_005|clock_xer|out_data_buffer[6]~q ),
	.src_data_6(src_data_6),
	.readdata_7(readdata_7),
	.av_readdata_pre_71(\adc_0_adc_slave_translator|av_readdata_pre[7]~q ),
	.readdata_71(readdata_71),
	.readdata_72(readdata_72),
	.out_data_buffer_7(\crosser_004|clock_xer|out_data_buffer[7]~q ),
	.readdata_73(readdata_73),
	.av_readdata_pre_72(\timer_0_s1_translator|av_readdata_pre[7]~q ),
	.out_data_buffer_71(\crosser_005|clock_xer|out_data_buffer[7]~q ),
	.src_data_7(src_data_7),
	.src_payload(src_payload10),
	.readdata_232(readdata_232),
	.out_data_buffer_23(\crosser_005|clock_xer|out_data_buffer[23]~q ),
	.src_payload1(src_payload11),
	.readdata_222(readdata_222),
	.out_data_buffer_22(\crosser_005|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_221(\crosser_004|clock_xer|out_data_buffer[22]~q ),
	.src_payload2(src_payload12),
	.readdata_212(readdata_213),
	.out_data_buffer_211(\crosser_005|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_212(\crosser_004|clock_xer|out_data_buffer[21]~q ),
	.src_payload3(src_payload13),
	.readdata_202(readdata_202),
	.out_data_buffer_20(\crosser_005|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_201(\crosser_004|clock_xer|out_data_buffer[20]~q ),
	.src_payload4(src_payload14),
	.readdata_192(readdata_192),
	.out_data_buffer_19(\crosser_005|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_191(\crosser_004|clock_xer|out_data_buffer[19]~q ),
	.src_payload5(src_payload15),
	.readdata_182(readdata_182),
	.out_data_buffer_18(\crosser_005|clock_xer|out_data_buffer[18]~q ),
	.out_data_buffer_181(\crosser_004|clock_xer|out_data_buffer[18]~q ),
	.src_payload6(src_payload16),
	.readdata_172(readdata_172),
	.out_data_buffer_17(\crosser_005|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_171(\crosser_004|clock_xer|out_data_buffer[17]~q ),
	.src_payload7(src_payload17),
	.readdata_162(readdata_163),
	.out_data_buffer_16(\crosser_005|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_161(\crosser_004|clock_xer|out_data_buffer[16]~q ),
	.src_payload8(src_payload18),
	.readdata_151(readdata_152),
	.av_readdata_pre_151(\adc_0_adc_slave_translator|av_readdata_pre[15]~q ),
	.readdata_152(readdata_153),
	.readdata_153(readdata_154),
	.out_data_buffer_15(\crosser_004|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_151(\crosser_005|clock_xer|out_data_buffer[15]~q ),
	.av_readdata_pre_152(\timer_0_s1_translator|av_readdata_pre[15]~q ),
	.src_data_151(src_data_151),
	.out_data_buffer_14(\crosser_004|clock_xer|out_data_buffer[14]~q ),
	.readdata_141(readdata_142),
	.av_readdata_pre_141(\timer_0_s1_translator|av_readdata_pre[14]~q ),
	.out_data_buffer_141(\crosser_005|clock_xer|out_data_buffer[14]~q ),
	.src_data_14(src_data_14),
	.av_readdata_pre_131(\timer_0_s1_translator|av_readdata_pre[13]~q ),
	.readdata_131(readdata_132),
	.out_data_buffer_13(\crosser_005|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_131(\crosser_004|clock_xer|out_data_buffer[13]~q ),
	.src_data_131(src_data_131),
	.out_data_buffer_121(\crosser_004|clock_xer|out_data_buffer[12]~q ),
	.readdata_121(readdata_122),
	.av_readdata_pre_121(\timer_0_s1_translator|av_readdata_pre[12]~q ),
	.out_data_buffer_122(\crosser_005|clock_xer|out_data_buffer[12]~q ),
	.src_data_121(src_data_121),
	.readdata_111(readdata_112),
	.av_readdata_pre_112(\adc_0_adc_slave_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_113(\timer_0_s1_translator|av_readdata_pre[11]~q ),
	.out_data_buffer_111(\crosser_005|clock_xer|out_data_buffer[11]~q ),
	.src_data_111(src_data_111),
	.av_readdata_pre_101(\timer_0_s1_translator|av_readdata_pre[10]~q ),
	.readdata_10(readdata_101),
	.av_readdata_pre_102(\adc_0_adc_slave_translator|av_readdata_pre[10]~q ),
	.out_data_buffer_10(\crosser_005|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_101(\crosser_004|clock_xer|out_data_buffer[10]~q ),
	.src_data_10(src_data_10),
	.readdata_9(readdata_91),
	.av_readdata_pre_91(\adc_0_adc_slave_translator|av_readdata_pre[9]~q ),
	.readdata_91(readdata_92),
	.readdata_92(readdata_93),
	.out_data_buffer_9(\crosser_004|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_91(\crosser_005|clock_xer|out_data_buffer[9]~q ),
	.av_readdata_pre_92(\timer_0_s1_translator|av_readdata_pre[9]~q ),
	.src_data_9(src_data_9),
	.readdata_8(readdata_81),
	.av_readdata_pre_81(\adc_0_adc_slave_translator|av_readdata_pre[8]~q ),
	.readdata_81(readdata_82),
	.readdata_82(readdata_83),
	.out_data_buffer_8(\crosser_004|clock_xer|out_data_buffer[8]~q ),
	.av_readdata_pre_82(\timer_0_s1_translator|av_readdata_pre[8]~q ),
	.out_data_buffer_81(\crosser_005|clock_xer|out_data_buffer[8]~q ),
	.src_data_8(src_data_8));

niosII_niosII_mm_interconnect_0_rsp_demux_009_2 rsp_demux_012(
	.rp_valid(\sdram_s1_agent|rp_valid~combout ),
	.always10(\sdram_s1_rsp_width_adapter|always10~1_combout ),
	.mem_66_0(\sdram_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_48_0(\sdram_s1_agent_rsp_fifo|mem[0][48]~q ),
	.src0_valid(src0_valid),
	.src1_valid(src1_valid1));

niosII_niosII_mm_interconnect_0_rsp_demux_009_1 rsp_demux_010(
	.mem_84_0(\epcs_epcs_control_port_agent_rsp_fifo|mem[0][84]~q ),
	.mem_66_0(\epcs_epcs_control_port_agent_rsp_fifo|mem[0][66]~q ),
	.in_data_toggle(\crosser_006|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser_006|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.in_data_toggle1(\crosser_005|clock_xer|in_data_toggle~q ),
	.dreg_01(\crosser_005|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.take_in_data(\crosser_006|clock_xer|take_in_data~0_combout ),
	.WideOr0(\rsp_demux_010|WideOr0~1_combout ));

niosII_niosII_mm_interconnect_0_rsp_demux_009 rsp_demux_009(
	.mem_84_0(mem_84_0),
	.mem_66_0(mem_66_0),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.src1_valid(src1_valid),
	.src0_valid(\rsp_demux_009|src0_valid~0_combout ));

niosII_niosII_mm_interconnect_0_cmd_mux_009_2 cmd_mux_012(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.r_sync_rst(r_sync_rst),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.cp_valid(cp_valid),
	.saved_grant_0(saved_grant_01),
	.saved_grant_1(saved_grant_11),
	.WideOr0(WideOr0),
	.Equal0(Equal0),
	.src_channel_12(\router|src_channel[12]~0_combout ),
	.src_channel_121(\router|src_channel[12]~3_combout ),
	.cp_valid1(\cpu_instruction_master_agent|cp_valid~combout ),
	.F_pc_22(F_pc_22),
	.F_pc_21(F_pc_21),
	.F_pc_20(F_pc_20),
	.F_pc_19(F_pc_19),
	.F_pc_18(F_pc_18),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.F_pc_10(F_pc_10),
	.Equal1(\router_001|Equal1~4_combout ),
	.Equal11(Equal1),
	.src_channel_122(\router|src_channel[12]~4_combout ),
	.WideOr11(WideOr1),
	.mem_used_7(mem_used_7),
	.uav_read1(\cpu_instruction_master_translator|uav_read~combout ),
	.src_data_66(src_data_66),
	.F_pc_8(F_pc_8),
	.src_data_46(\cmd_mux_012|src_data[46]~combout ),
	.src_valid(src_valid2),
	.src_data_60(\cmd_mux_012|src_data[60]~combout ),
	.F_pc_9(F_pc_9),
	.src_data_47(\cmd_mux_012|src_data[47]~combout ),
	.src_data_49(\cmd_mux_012|src_data[49]~combout ),
	.src_data_48(\cmd_mux_012|src_data[48]~combout ),
	.src_data_51(\cmd_mux_012|src_data[51]~combout ),
	.src_data_50(\cmd_mux_012|src_data[50]~combout ),
	.src_data_53(\cmd_mux_012|src_data[53]~combout ),
	.src_data_52(\cmd_mux_012|src_data[52]~combout ),
	.src_data_55(\cmd_mux_012|src_data[55]~combout ),
	.src_data_54(\cmd_mux_012|src_data[54]~combout ),
	.src_data_57(\cmd_mux_012|src_data[57]~combout ),
	.src_data_56(\cmd_mux_012|src_data[56]~combout ),
	.src_data_59(\cmd_mux_012|src_data[59]~combout ),
	.src_data_58(\cmd_mux_012|src_data[58]~combout ),
	.F_pc_0(F_pc_0),
	.src_data_38(\cmd_mux_012|src_data[38]~combout ),
	.F_pc_1(F_pc_1),
	.src_data_39(\cmd_mux_012|src_data[39]~combout ),
	.F_pc_2(F_pc_2),
	.src_data_40(\cmd_mux_012|src_data[40]~combout ),
	.F_pc_3(F_pc_3),
	.src_data_41(\cmd_mux_012|src_data[41]~combout ),
	.F_pc_4(F_pc_4),
	.src_data_42(\cmd_mux_012|src_data[42]~combout ),
	.F_pc_5(F_pc_5),
	.src_data_43(\cmd_mux_012|src_data[43]~combout ),
	.F_pc_6(F_pc_6),
	.src_data_44(\cmd_mux_012|src_data[44]~combout ),
	.F_pc_7(F_pc_7),
	.src_data_45(\cmd_mux_012|src_data[45]~combout ),
	.count_0(\sdram_s1_cmd_width_adapter|count[0]~q ),
	.last_cycle(\cmd_mux_012|last_cycle~0_combout ),
	.src12_valid(\cmd_demux|src12_valid~2_combout ),
	.src_payload_0(\cmd_mux_012|src_payload[0]~combout ),
	.d_byteenable_2(d_byteenable_2),
	.src_data_34(\cmd_mux_012|src_data[34]~combout ),
	.d_byteenable_3(d_byteenable_3),
	.src_data_35(\cmd_mux_012|src_data[35]~combout ),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.src_payload(\cmd_mux_012|src_payload~0_combout ),
	.src_payload1(\cmd_mux_012|src_payload~1_combout ),
	.src_payload2(\cmd_mux_012|src_payload~2_combout ),
	.src_payload3(\cmd_mux_012|src_payload~3_combout ),
	.src_payload4(\cmd_mux_012|src_payload~4_combout ),
	.src_payload5(\cmd_mux_012|src_payload~5_combout ),
	.src_payload6(\cmd_mux_012|src_payload~6_combout ),
	.src_payload7(\cmd_mux_012|src_payload~7_combout ),
	.src_payload8(\cmd_mux_012|src_payload~8_combout ),
	.src_payload9(\cmd_mux_012|src_payload~9_combout ),
	.src_payload10(\cmd_mux_012|src_payload~10_combout ),
	.src_payload11(\cmd_mux_012|src_payload~11_combout ),
	.src_payload12(\cmd_mux_012|src_payload~12_combout ),
	.src_payload13(\cmd_mux_012|src_payload~13_combout ),
	.src_payload14(\cmd_mux_012|src_payload~14_combout ),
	.src_payload15(\cmd_mux_012|src_payload~15_combout ),
	.src2_valid(\cmd_demux_001|src2_valid~2_combout ));

niosII_niosII_mm_interconnect_0_cmd_mux_009_1 cmd_mux_010(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst1),
	.saved_grant_0(saved_grant_0),
	.saved_grant_1(saved_grant_1),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_381(\crosser_001|clock_xer|out_data_buffer[38]~q ),
	.src_data_38(src_data_38),
	.out_data_buffer_39(\crosser_003|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_391(\crosser_001|clock_xer|out_data_buffer[39]~q ),
	.src_data_39(src_data_39),
	.out_data_buffer_40(\crosser_003|clock_xer|out_data_buffer[40]~q ),
	.out_data_buffer_401(\crosser_001|clock_xer|out_data_buffer[40]~q ),
	.src_data_40(src_data_40),
	.out_data_buffer_10(\crosser_001|clock_xer|out_data_buffer[10]~q ),
	.src_payload(src_payload),
	.out_data_buffer_0(\crosser_001|clock_xer|out_data_buffer[0]~q ),
	.src_payload1(src_payload1),
	.out_data_toggle_flopped(\crosser_001|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_001|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(\crosser_001|clock_xer|out_valid~combout ),
	.out_data_toggle_flopped1(\crosser_003|clock_xer|out_data_toggle_flopped~q ),
	.dreg_01(\crosser_003|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid1(\crosser_003|clock_xer|out_valid~combout ),
	.wait_latency_counter_0(\epcs_epcs_control_port_translator|wait_latency_counter[0]~q ),
	.waitrequest_reset_override(\epcs_epcs_control_port_translator|waitrequest_reset_override~q ),
	.mem_used_1(mem_used_11),
	.wait_latency_counter_1(wait_latency_counter_1),
	.last_cycle(\cmd_mux_010|last_cycle~0_combout ),
	.out_data_buffer_105(\crosser_003|clock_xer|out_data_buffer[105]~q ),
	.out_data_buffer_1051(\crosser_001|clock_xer|out_data_buffer[105]~q ),
	.src_payload_0(\cmd_mux_010|src_payload[0]~combout ),
	.src_valid(src_valid),
	.src_valid1(src_valid1),
	.out_data_buffer_46(\crosser_003|clock_xer|out_data_buffer[46]~q ),
	.out_data_buffer_461(\crosser_001|clock_xer|out_data_buffer[46]~q ),
	.src_data_46(src_data_46),
	.out_data_buffer_7(\crosser_001|clock_xer|out_data_buffer[7]~q ),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.out_data_buffer_66(\crosser_003|clock_xer|out_data_buffer[66]~q ),
	.out_data_buffer_661(\crosser_001|clock_xer|out_data_buffer[66]~q ),
	.src_data_66(src_data_661),
	.out_data_buffer_6(\crosser_001|clock_xer|out_data_buffer[6]~q ),
	.src_payload4(src_payload4),
	.out_data_buffer_5(\crosser_001|clock_xer|out_data_buffer[5]~q ),
	.src_payload5(src_payload5),
	.out_data_buffer_4(\crosser_001|clock_xer|out_data_buffer[4]~q ),
	.src_payload6(src_payload7),
	.out_data_buffer_3(\crosser_001|clock_xer|out_data_buffer[3]~q ),
	.src_payload7(src_payload19),
	.out_data_buffer_2(\crosser_001|clock_xer|out_data_buffer[2]~q ),
	.src_payload8(src_payload21),
	.out_data_buffer_1(\crosser_001|clock_xer|out_data_buffer[1]~q ),
	.src_payload9(src_payload25),
	.out_data_buffer_41(\crosser_003|clock_xer|out_data_buffer[41]~q ),
	.out_data_buffer_411(\crosser_001|clock_xer|out_data_buffer[41]~q ),
	.src_data_41(src_data_412),
	.out_data_buffer_42(\crosser_003|clock_xer|out_data_buffer[42]~q ),
	.out_data_buffer_421(\crosser_001|clock_xer|out_data_buffer[42]~q ),
	.src_data_42(src_data_421),
	.out_data_buffer_43(\crosser_003|clock_xer|out_data_buffer[43]~q ),
	.out_data_buffer_431(\crosser_001|clock_xer|out_data_buffer[43]~q ),
	.src_data_43(src_data_431),
	.out_data_buffer_44(\crosser_003|clock_xer|out_data_buffer[44]~q ),
	.out_data_buffer_441(\crosser_001|clock_xer|out_data_buffer[44]~q ),
	.src_data_44(src_data_441),
	.out_data_buffer_45(\crosser_003|clock_xer|out_data_buffer[45]~q ),
	.out_data_buffer_451(\crosser_001|clock_xer|out_data_buffer[45]~q ),
	.src_data_45(src_data_451),
	.src_payload10(src_payload26),
	.out_data_buffer_11(\crosser_001|clock_xer|out_data_buffer[11]~q ),
	.src_payload11(src_payload53),
	.out_data_buffer_13(\crosser_001|clock_xer|out_data_buffer[13]~q ),
	.src_payload12(src_payload54),
	.out_data_buffer_12(\crosser_001|clock_xer|out_data_buffer[12]~q ),
	.src_payload13(src_payload55),
	.out_data_buffer_14(\crosser_001|clock_xer|out_data_buffer[14]~q ),
	.src_payload14(src_payload56),
	.out_data_buffer_15(\crosser_001|clock_xer|out_data_buffer[15]~q ),
	.src_payload15(src_payload57),
	.out_data_buffer_9(\crosser_001|clock_xer|out_data_buffer[9]~q ),
	.src_payload16(src_payload59),
	.out_data_buffer_8(\crosser_001|clock_xer|out_data_buffer[8]~q ),
	.src_payload17(src_payload60),
	.WideOr11(\cmd_mux_010|WideOr1~combout ));

niosII_niosII_mm_interconnect_0_cmd_mux_009 cmd_mux_009(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.r_sync_rst(r_sync_rst),
	.cp_valid(cp_valid),
	.d_writedata_0(d_writedata_0),
	.d_byteenable_0(d_byteenable_0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_byteenable_1(d_byteenable_1),
	.Equal2(\router|Equal2~1_combout ),
	.F_pc_8(F_pc_8),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.F_pc_2(F_pc_2),
	.F_pc_3(F_pc_3),
	.F_pc_4(F_pc_4),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_7(F_pc_7),
	.saved_grant_0(saved_grant_02),
	.waitrequest(waitrequest1),
	.mem_used_1(mem_used_15),
	.d_writedata_10(d_writedata_10),
	.d_byteenable_2(d_byteenable_2),
	.d_byteenable_3(d_byteenable_3),
	.saved_grant_1(\cmd_mux_009|saved_grant[1]~q ),
	.hbreak_enabled(hbreak_enabled),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.WideOr11(WideOr12),
	.src_data_46(src_data_461),
	.src_payload(src_payload8),
	.src_payload1(src_payload9),
	.src_data_38(src_data_381),
	.src_data_39(src_data_391),
	.src_data_40(src_data_401),
	.src_data_41(src_data_411),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_32(src_data_32),
	.src_payload2(src_payload20),
	.src_payload3(src_payload22),
	.src_payload4(src_payload23),
	.src_payload5(src_payload24),
	.src_payload6(src_payload27),
	.src_data_33(src_data_33),
	.src_payload7(src_payload28),
	.src_payload8(src_payload29),
	.src_data_34(src_data_34),
	.src_payload9(src_payload30),
	.src_payload10(src_payload31),
	.src_payload11(src_payload32),
	.src_payload12(src_payload33),
	.src_payload13(src_payload34),
	.src_payload14(src_payload35),
	.src_payload15(src_payload36),
	.src_payload16(src_payload37),
	.src_payload17(src_payload38),
	.src_payload18(src_payload39),
	.src_payload19(src_payload40),
	.src_data_35(src_data_35),
	.src_payload20(src_payload41),
	.src_payload21(src_payload42),
	.src_payload22(src_payload43),
	.src_payload23(src_payload44),
	.src_payload24(src_payload45),
	.src_payload25(src_payload46),
	.src_payload26(src_payload47),
	.src_payload27(src_payload48),
	.src_payload28(src_payload49),
	.src_payload29(src_payload50),
	.src_payload30(src_payload51),
	.src_payload31(src_payload52),
	.src_payload32(src_payload58));

niosII_altera_avalon_st_handshake_clock_crosser_7 crosser_007(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.out_data_toggle_flopped(\crosser_007|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_007|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.in_ready(\crosser_007|clock_xer|in_ready~0_combout ),
	.rp_valid(\sys_pll_pll_slave_agent|rp_valid~combout ),
	.out_valid(\crosser_007|clock_xer|out_valid~combout ),
	.out_data_buffer_0(\crosser_007|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_1(\crosser_007|clock_xer|out_data_buffer[1]~q ),
	.out_data_0(\sys_pll_pll_slave_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\sys_pll_pll_slave_agent_rdata_fifo|out_data[1]~1_combout ),
	.clk_clk(clk_clk));

niosII_altera_avalon_st_handshake_clock_crosser_6 crosser_006(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.r_sync_rst1(r_sync_rst1),
	.mem_84_0(\epcs_epcs_control_port_agent_rsp_fifo|mem[0][84]~q ),
	.mem_66_0(\epcs_epcs_control_port_agent_rsp_fifo|mem[0][66]~q ),
	.in_data_toggle(\crosser_006|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser_006|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.take_in_data(\crosser_006|clock_xer|take_in_data~0_combout ),
	.out_data_toggle_flopped(\crosser_006|clock_xer|out_data_toggle_flopped~q ),
	.dreg_01(\crosser_006|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.rp_valid(\epcs_epcs_control_port_agent|rp_valid~combout ),
	.out_valid(out_valid),
	.out_data_buffer_0(out_data_buffer_01),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_0(\epcs_epcs_control_port_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\epcs_epcs_control_port_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\epcs_epcs_control_port_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\epcs_epcs_control_port_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\epcs_epcs_control_port_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_11(\epcs_epcs_control_port_agent_rdata_fifo|out_data[11]~5_combout ),
	.out_data_13(\epcs_epcs_control_port_agent_rdata_fifo|out_data[13]~6_combout ),
	.out_data_16(\epcs_epcs_control_port_agent_rdata_fifo|out_data[16]~7_combout ),
	.out_data_12(\epcs_epcs_control_port_agent_rdata_fifo|out_data[12]~8_combout ),
	.out_data_5(\epcs_epcs_control_port_agent_rdata_fifo|out_data[5]~9_combout ),
	.out_data_14(\epcs_epcs_control_port_agent_rdata_fifo|out_data[14]~10_combout ),
	.out_data_15(\epcs_epcs_control_port_agent_rdata_fifo|out_data[15]~11_combout ),
	.out_data_10(\epcs_epcs_control_port_agent_rdata_fifo|out_data[10]~12_combout ),
	.out_data_9(\epcs_epcs_control_port_agent_rdata_fifo|out_data[9]~13_combout ),
	.out_data_8(\epcs_epcs_control_port_agent_rdata_fifo|out_data[8]~14_combout ),
	.out_data_7(\epcs_epcs_control_port_agent_rdata_fifo|out_data[7]~15_combout ),
	.out_data_6(\epcs_epcs_control_port_agent_rdata_fifo|out_data[6]~16_combout ),
	.out_data_21(\epcs_epcs_control_port_agent_rdata_fifo|out_data[21]~17_combout ),
	.out_data_30(\epcs_epcs_control_port_agent_rdata_fifo|out_data[30]~18_combout ),
	.out_data_29(\epcs_epcs_control_port_agent_rdata_fifo|out_data[29]~19_combout ),
	.out_data_28(\epcs_epcs_control_port_agent_rdata_fifo|out_data[28]~20_combout ),
	.out_data_27(\epcs_epcs_control_port_agent_rdata_fifo|out_data[27]~21_combout ),
	.out_data_26(\epcs_epcs_control_port_agent_rdata_fifo|out_data[26]~22_combout ),
	.out_data_25(\epcs_epcs_control_port_agent_rdata_fifo|out_data[25]~23_combout ),
	.out_data_24(\epcs_epcs_control_port_agent_rdata_fifo|out_data[24]~24_combout ),
	.out_data_23(\epcs_epcs_control_port_agent_rdata_fifo|out_data[23]~25_combout ),
	.out_data_22(\epcs_epcs_control_port_agent_rdata_fifo|out_data[22]~26_combout ),
	.out_data_20(\epcs_epcs_control_port_agent_rdata_fifo|out_data[20]~27_combout ),
	.out_data_19(\epcs_epcs_control_port_agent_rdata_fifo|out_data[19]~28_combout ),
	.out_data_18(\epcs_epcs_control_port_agent_rdata_fifo|out_data[18]~29_combout ),
	.out_data_17(\epcs_epcs_control_port_agent_rdata_fifo|out_data[17]~30_combout ),
	.out_data_31(\epcs_epcs_control_port_agent_rdata_fifo|out_data[31]~31_combout ));

endmodule

module niosII_altera_avalon_sc_fifo (
	clk,
	reset,
	mem_used_1,
	uav_read,
	hold_waitrequest,
	Equal3,
	read_latency_shift_reg_0,
	waitrequest,
	m0_read,
	read_latency_shift_reg)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
output 	mem_used_1;
input 	uav_read;
input 	hold_waitrequest;
input 	Equal3;
input 	read_latency_shift_reg_0;
input 	waitrequest;
input 	m0_read;
input 	read_latency_shift_reg;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~2_combout ),
	.datab(m0_read),
	.datac(read_latency_shift_reg),
	.datad(waitrequest),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(hold_waitrequest),
	.datab(uav_read),
	.datac(Equal3),
	.datad(waitrequest),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_1 (
	clk,
	reset,
	uav_read,
	uav_read1,
	mem_84_0,
	mem_66_0,
	read_latency_shift_reg_0,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	write,
	saved_grant_1,
	mem,
	WideOr1,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	uav_read;
input 	uav_read1;
output 	mem_84_0;
output 	mem_66_0;
input 	read_latency_shift_reg_0;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
output 	write;
input 	saved_grant_1;
output 	mem;
input 	WideOr1;
input 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][84]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][66]~q ;
wire \mem~2_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][84] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_84_0),
	.prn(vcc));
defparam \mem[0][84] .is_wysiwyg = "true";
defparam \mem[0][84] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(write),
	.cout());
defparam \write~0 .lut_mask = 16'h0FFF;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~1 (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(mem),
	.cout());
defparam \mem~1 .lut_mask = 16'hFFFE;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][84] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][84]~q ),
	.prn(vcc));
defparam \mem[1][84] .is_wysiwyg = "true";
defparam \mem[1][84] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][84]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(write),
	.datac(WideOr1),
	.datad(mem),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][66]~q ),
	.datab(mem),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hAFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(rf_source_valid),
	.datac(\mem_used[1]~0_combout ),
	.datad(waitrequest),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_2 (
	clk,
	reset,
	mem_used_0,
	mem_105_0,
	read_latency_shift_reg_0,
	mem_used_01,
	rp_valid,
	WideOr0,
	av_readdata_pre_0,
	out_data_0,
	av_readdata_pre_1,
	out_data_1,
	av_readdata_pre_2,
	out_data_2,
	av_readdata_pre_3,
	out_data_3,
	av_readdata_pre_4,
	out_data_4,
	av_readdata_pre_11,
	out_data_11,
	av_readdata_pre_13,
	out_data_13,
	av_readdata_pre_16,
	out_data_16,
	av_readdata_pre_12,
	out_data_12,
	av_readdata_pre_5,
	out_data_5,
	av_readdata_pre_14,
	out_data_14,
	av_readdata_pre_15,
	out_data_15,
	av_readdata_pre_10,
	out_data_10,
	av_readdata_pre_9,
	out_data_9,
	av_readdata_pre_8,
	out_data_8,
	av_readdata_pre_7,
	out_data_7,
	av_readdata_pre_6,
	out_data_6,
	av_readdata_pre_21,
	out_data_21,
	av_readdata_pre_30,
	out_data_30,
	av_readdata_pre_29,
	out_data_29,
	av_readdata_pre_28,
	out_data_28,
	av_readdata_pre_27,
	out_data_27,
	av_readdata_pre_26,
	out_data_26,
	av_readdata_pre_25,
	out_data_25,
	av_readdata_pre_24,
	out_data_24,
	av_readdata_pre_23,
	out_data_23,
	av_readdata_pre_22,
	out_data_22,
	av_readdata_pre_20,
	out_data_20,
	av_readdata_pre_19,
	out_data_19,
	av_readdata_pre_18,
	out_data_18,
	av_readdata_pre_17,
	out_data_17,
	av_readdata_pre_31,
	out_data_31)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	mem_used_0;
input 	mem_105_0;
input 	read_latency_shift_reg_0;
output 	mem_used_01;
input 	rp_valid;
input 	WideOr0;
input 	av_readdata_pre_0;
output 	out_data_0;
input 	av_readdata_pre_1;
output 	out_data_1;
input 	av_readdata_pre_2;
output 	out_data_2;
input 	av_readdata_pre_3;
output 	out_data_3;
input 	av_readdata_pre_4;
output 	out_data_4;
input 	av_readdata_pre_11;
output 	out_data_11;
input 	av_readdata_pre_13;
output 	out_data_13;
input 	av_readdata_pre_16;
output 	out_data_16;
input 	av_readdata_pre_12;
output 	out_data_12;
input 	av_readdata_pre_5;
output 	out_data_5;
input 	av_readdata_pre_14;
output 	out_data_14;
input 	av_readdata_pre_15;
output 	out_data_15;
input 	av_readdata_pre_10;
output 	out_data_10;
input 	av_readdata_pre_9;
output 	out_data_9;
input 	av_readdata_pre_8;
output 	out_data_8;
input 	av_readdata_pre_7;
output 	out_data_7;
input 	av_readdata_pre_6;
output 	out_data_6;
input 	av_readdata_pre_21;
output 	out_data_21;
input 	av_readdata_pre_30;
output 	out_data_30;
input 	av_readdata_pre_29;
output 	out_data_29;
input 	av_readdata_pre_28;
output 	out_data_28;
input 	av_readdata_pre_27;
output 	out_data_27;
input 	av_readdata_pre_26;
output 	out_data_26;
input 	av_readdata_pre_25;
output 	out_data_25;
input 	av_readdata_pre_24;
output 	out_data_24;
input 	av_readdata_pre_23;
output 	out_data_23;
input 	av_readdata_pre_22;
output 	out_data_22;
input 	av_readdata_pre_20;
output 	out_data_20;
input 	av_readdata_pre_19;
output 	out_data_19;
input 	av_readdata_pre_18;
output 	out_data_18;
input 	av_readdata_pre_17;
output 	out_data_17;
input 	av_readdata_pre_31;
output 	out_data_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~4_combout ;
wire \mem[0][0]~q ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[0][1]~q ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[0][2]~q ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[0][3]~q ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[0][4]~q ;
wire \mem[1][11]~q ;
wire \mem~5_combout ;
wire \mem[0][11]~q ;
wire \mem[1][13]~q ;
wire \mem~6_combout ;
wire \mem[0][13]~q ;
wire \mem[1][16]~q ;
wire \mem~7_combout ;
wire \mem[0][16]~q ;
wire \mem[1][12]~q ;
wire \mem~8_combout ;
wire \mem[0][12]~q ;
wire \mem[1][5]~q ;
wire \mem~9_combout ;
wire \mem[0][5]~q ;
wire \mem[1][14]~q ;
wire \mem~10_combout ;
wire \mem[0][14]~q ;
wire \mem[1][15]~q ;
wire \mem~11_combout ;
wire \mem[0][15]~q ;
wire \mem[1][10]~q ;
wire \mem~12_combout ;
wire \mem[0][10]~q ;
wire \mem[1][9]~q ;
wire \mem~13_combout ;
wire \mem[0][9]~q ;
wire \mem[1][8]~q ;
wire \mem~14_combout ;
wire \mem[0][8]~q ;
wire \mem[1][7]~q ;
wire \mem~15_combout ;
wire \mem[0][7]~q ;
wire \mem[1][6]~q ;
wire \mem~16_combout ;
wire \mem[0][6]~q ;
wire \mem[1][21]~q ;
wire \mem~17_combout ;
wire \mem[0][21]~q ;
wire \mem[1][30]~q ;
wire \mem~18_combout ;
wire \mem[0][30]~q ;
wire \mem[1][29]~q ;
wire \mem~19_combout ;
wire \mem[0][29]~q ;
wire \mem[1][28]~q ;
wire \mem~20_combout ;
wire \mem[0][28]~q ;
wire \mem[1][27]~q ;
wire \mem~21_combout ;
wire \mem[0][27]~q ;
wire \mem[1][26]~q ;
wire \mem~22_combout ;
wire \mem[0][26]~q ;
wire \mem[1][25]~q ;
wire \mem~23_combout ;
wire \mem[0][25]~q ;
wire \mem[1][24]~q ;
wire \mem~24_combout ;
wire \mem[0][24]~q ;
wire \mem[1][23]~q ;
wire \mem~25_combout ;
wire \mem[0][23]~q ;
wire \mem[1][22]~q ;
wire \mem~26_combout ;
wire \mem[0][22]~q ;
wire \mem[1][20]~q ;
wire \mem~27_combout ;
wire \mem[0][20]~q ;
wire \mem[1][19]~q ;
wire \mem~28_combout ;
wire \mem[0][19]~q ;
wire \mem[1][18]~q ;
wire \mem~29_combout ;
wire \mem[0][18]~q ;
wire \mem[1][17]~q ;
wire \mem~30_combout ;
wire \mem[0][17]~q ;
wire \mem[1][31]~q ;
wire \mem~31_combout ;
wire \mem[0][31]~q ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_01),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \out_data[0]~0 (
	.dataa(\mem[0][0]~q ),
	.datab(av_readdata_pre_0),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_0),
	.cout());
defparam \out_data[0]~0 .lut_mask = 16'hEFFE;
defparam \out_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[1]~1 (
	.dataa(\mem[0][1]~q ),
	.datab(av_readdata_pre_1),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_1),
	.cout());
defparam \out_data[1]~1 .lut_mask = 16'hEFFE;
defparam \out_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[2]~2 (
	.dataa(\mem[0][2]~q ),
	.datab(av_readdata_pre_2),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_2),
	.cout());
defparam \out_data[2]~2 .lut_mask = 16'hEFFE;
defparam \out_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[3]~3 (
	.dataa(\mem[0][3]~q ),
	.datab(av_readdata_pre_3),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_3),
	.cout());
defparam \out_data[3]~3 .lut_mask = 16'hEFFE;
defparam \out_data[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[4]~4 (
	.dataa(\mem[0][4]~q ),
	.datab(av_readdata_pre_4),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_4),
	.cout());
defparam \out_data[4]~4 .lut_mask = 16'hEFFE;
defparam \out_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[11]~5 (
	.dataa(\mem[0][11]~q ),
	.datab(av_readdata_pre_11),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_11),
	.cout());
defparam \out_data[11]~5 .lut_mask = 16'hEFFE;
defparam \out_data[11]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[13]~6 (
	.dataa(\mem[0][13]~q ),
	.datab(av_readdata_pre_13),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_13),
	.cout());
defparam \out_data[13]~6 .lut_mask = 16'hEFFE;
defparam \out_data[13]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[16]~7 (
	.dataa(\mem[0][16]~q ),
	.datab(av_readdata_pre_16),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_16),
	.cout());
defparam \out_data[16]~7 .lut_mask = 16'hEFFE;
defparam \out_data[16]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[12]~8 (
	.dataa(\mem[0][12]~q ),
	.datab(av_readdata_pre_12),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_12),
	.cout());
defparam \out_data[12]~8 .lut_mask = 16'hEFFE;
defparam \out_data[12]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[5]~9 (
	.dataa(\mem[0][5]~q ),
	.datab(av_readdata_pre_5),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_5),
	.cout());
defparam \out_data[5]~9 .lut_mask = 16'hEFFE;
defparam \out_data[5]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[14]~10 (
	.dataa(\mem[0][14]~q ),
	.datab(av_readdata_pre_14),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_14),
	.cout());
defparam \out_data[14]~10 .lut_mask = 16'hEFFE;
defparam \out_data[14]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[15]~11 (
	.dataa(\mem[0][15]~q ),
	.datab(av_readdata_pre_15),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_15),
	.cout());
defparam \out_data[15]~11 .lut_mask = 16'hEFFE;
defparam \out_data[15]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[10]~12 (
	.dataa(\mem[0][10]~q ),
	.datab(av_readdata_pre_10),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_10),
	.cout());
defparam \out_data[10]~12 .lut_mask = 16'hEFFE;
defparam \out_data[10]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[9]~13 (
	.dataa(\mem[0][9]~q ),
	.datab(av_readdata_pre_9),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_9),
	.cout());
defparam \out_data[9]~13 .lut_mask = 16'hEFFE;
defparam \out_data[9]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[8]~14 (
	.dataa(\mem[0][8]~q ),
	.datab(av_readdata_pre_8),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_8),
	.cout());
defparam \out_data[8]~14 .lut_mask = 16'hEFFE;
defparam \out_data[8]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[7]~15 (
	.dataa(\mem[0][7]~q ),
	.datab(av_readdata_pre_7),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_7),
	.cout());
defparam \out_data[7]~15 .lut_mask = 16'hEFFE;
defparam \out_data[7]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[6]~16 (
	.dataa(\mem[0][6]~q ),
	.datab(av_readdata_pre_6),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_6),
	.cout());
defparam \out_data[6]~16 .lut_mask = 16'hEFFE;
defparam \out_data[6]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[21]~17 (
	.dataa(\mem[0][21]~q ),
	.datab(av_readdata_pre_21),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_21),
	.cout());
defparam \out_data[21]~17 .lut_mask = 16'hEFFE;
defparam \out_data[21]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[30]~18 (
	.dataa(\mem[0][30]~q ),
	.datab(av_readdata_pre_30),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_30),
	.cout());
defparam \out_data[30]~18 .lut_mask = 16'hEFFE;
defparam \out_data[30]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[29]~19 (
	.dataa(\mem[0][29]~q ),
	.datab(av_readdata_pre_29),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_29),
	.cout());
defparam \out_data[29]~19 .lut_mask = 16'hEFFE;
defparam \out_data[29]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[28]~20 (
	.dataa(\mem[0][28]~q ),
	.datab(av_readdata_pre_28),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_28),
	.cout());
defparam \out_data[28]~20 .lut_mask = 16'hEFFE;
defparam \out_data[28]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[27]~21 (
	.dataa(\mem[0][27]~q ),
	.datab(av_readdata_pre_27),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_27),
	.cout());
defparam \out_data[27]~21 .lut_mask = 16'hEFFE;
defparam \out_data[27]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[26]~22 (
	.dataa(\mem[0][26]~q ),
	.datab(av_readdata_pre_26),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_26),
	.cout());
defparam \out_data[26]~22 .lut_mask = 16'hEFFE;
defparam \out_data[26]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[25]~23 (
	.dataa(\mem[0][25]~q ),
	.datab(av_readdata_pre_25),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_25),
	.cout());
defparam \out_data[25]~23 .lut_mask = 16'hEFFE;
defparam \out_data[25]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[24]~24 (
	.dataa(\mem[0][24]~q ),
	.datab(av_readdata_pre_24),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_24),
	.cout());
defparam \out_data[24]~24 .lut_mask = 16'hEFFE;
defparam \out_data[24]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[23]~25 (
	.dataa(\mem[0][23]~q ),
	.datab(av_readdata_pre_23),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_23),
	.cout());
defparam \out_data[23]~25 .lut_mask = 16'hEFFE;
defparam \out_data[23]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[22]~26 (
	.dataa(\mem[0][22]~q ),
	.datab(av_readdata_pre_22),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_22),
	.cout());
defparam \out_data[22]~26 .lut_mask = 16'hEFFE;
defparam \out_data[22]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[20]~27 (
	.dataa(\mem[0][20]~q ),
	.datab(av_readdata_pre_20),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_20),
	.cout());
defparam \out_data[20]~27 .lut_mask = 16'hEFFE;
defparam \out_data[20]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[19]~28 (
	.dataa(\mem[0][19]~q ),
	.datab(av_readdata_pre_19),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_19),
	.cout());
defparam \out_data[19]~28 .lut_mask = 16'hEFFE;
defparam \out_data[19]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[18]~29 (
	.dataa(\mem[0][18]~q ),
	.datab(av_readdata_pre_18),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_18),
	.cout());
defparam \out_data[18]~29 .lut_mask = 16'hEFFE;
defparam \out_data[18]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[17]~30 (
	.dataa(\mem[0][17]~q ),
	.datab(av_readdata_pre_17),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_17),
	.cout());
defparam \out_data[17]~30 .lut_mask = 16'hEFFE;
defparam \out_data[17]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[31]~31 (
	.dataa(\mem[0][31]~q ),
	.datab(av_readdata_pre_31),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_31),
	.cout());
defparam \out_data[31]~31 .lut_mask = 16'hEFFE;
defparam \out_data[31]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(mem_used_0),
	.datab(mem_105_0),
	.datac(WideOr0),
	.datad(rp_valid),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h7FFF;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[1]~q ),
	.datab(read_latency_shift_reg_0),
	.datac(mem_used_01),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~0 (
	.dataa(\mem_used[1]~q ),
	.datab(mem_used_01),
	.datac(read_latency_shift_reg_0),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~0_combout ),
	.cout());
defparam \mem_used[0]~0 .lut_mask = 16'hFDFE;
defparam \mem_used[0]~0 .sum_lutc_input = "datac";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][0]~q ),
	.datab(av_readdata_pre_0),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~4 (
	.dataa(mem_used_0),
	.datab(mem_105_0),
	.datac(mem_used_01),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\always0~4_combout ),
	.cout());
defparam \always0~4 .lut_mask = 16'h7FFF;
defparam \always0~4 .sum_lutc_input = "datac";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][0]~q ),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][1]~q ),
	.datab(av_readdata_pre_1),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][1]~q ),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][2]~q ),
	.datab(av_readdata_pre_2),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][2]~q ),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][3]~q ),
	.datab(av_readdata_pre_3),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hAACC;
defparam \mem~3 .sum_lutc_input = "datac";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][3]~q ),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[1][4]~q ),
	.datab(av_readdata_pre_4),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hAACC;
defparam \mem~4 .sum_lutc_input = "datac";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][4]~q ),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cycloneive_lcell_comb \mem~5 (
	.dataa(\mem[1][11]~q ),
	.datab(av_readdata_pre_11),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~5_combout ),
	.cout());
defparam \mem~5 .lut_mask = 16'hAACC;
defparam \mem~5 .sum_lutc_input = "datac";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][11]~q ),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cycloneive_lcell_comb \mem~6 (
	.dataa(\mem[1][13]~q ),
	.datab(av_readdata_pre_13),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~6_combout ),
	.cout());
defparam \mem~6 .lut_mask = 16'hAACC;
defparam \mem~6 .sum_lutc_input = "datac";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][13]~q ),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cycloneive_lcell_comb \mem~7 (
	.dataa(\mem[1][16]~q ),
	.datab(av_readdata_pre_16),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~7_combout ),
	.cout());
defparam \mem~7 .lut_mask = 16'hAACC;
defparam \mem~7 .sum_lutc_input = "datac";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][16]~q ),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cycloneive_lcell_comb \mem~8 (
	.dataa(\mem[1][12]~q ),
	.datab(av_readdata_pre_12),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~8_combout ),
	.cout());
defparam \mem~8 .lut_mask = 16'hAACC;
defparam \mem~8 .sum_lutc_input = "datac";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][12]~q ),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cycloneive_lcell_comb \mem~9 (
	.dataa(\mem[1][5]~q ),
	.datab(av_readdata_pre_5),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~9_combout ),
	.cout());
defparam \mem~9 .lut_mask = 16'hAACC;
defparam \mem~9 .sum_lutc_input = "datac";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][5]~q ),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cycloneive_lcell_comb \mem~10 (
	.dataa(\mem[1][14]~q ),
	.datab(av_readdata_pre_14),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~10_combout ),
	.cout());
defparam \mem~10 .lut_mask = 16'hAACC;
defparam \mem~10 .sum_lutc_input = "datac";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][14]~q ),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cycloneive_lcell_comb \mem~11 (
	.dataa(\mem[1][15]~q ),
	.datab(av_readdata_pre_15),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~11_combout ),
	.cout());
defparam \mem~11 .lut_mask = 16'hAACC;
defparam \mem~11 .sum_lutc_input = "datac";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][15]~q ),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cycloneive_lcell_comb \mem~12 (
	.dataa(\mem[1][10]~q ),
	.datab(av_readdata_pre_10),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~12_combout ),
	.cout());
defparam \mem~12 .lut_mask = 16'hAACC;
defparam \mem~12 .sum_lutc_input = "datac";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][10]~q ),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cycloneive_lcell_comb \mem~13 (
	.dataa(\mem[1][9]~q ),
	.datab(av_readdata_pre_9),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~13_combout ),
	.cout());
defparam \mem~13 .lut_mask = 16'hAACC;
defparam \mem~13 .sum_lutc_input = "datac";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][9]~q ),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cycloneive_lcell_comb \mem~14 (
	.dataa(\mem[1][8]~q ),
	.datab(av_readdata_pre_8),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~14_combout ),
	.cout());
defparam \mem~14 .lut_mask = 16'hAACC;
defparam \mem~14 .sum_lutc_input = "datac";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][8]~q ),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cycloneive_lcell_comb \mem~15 (
	.dataa(\mem[1][7]~q ),
	.datab(av_readdata_pre_7),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~15_combout ),
	.cout());
defparam \mem~15 .lut_mask = 16'hAACC;
defparam \mem~15 .sum_lutc_input = "datac";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][7]~q ),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cycloneive_lcell_comb \mem~16 (
	.dataa(\mem[1][6]~q ),
	.datab(av_readdata_pre_6),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~16_combout ),
	.cout());
defparam \mem~16 .lut_mask = 16'hAACC;
defparam \mem~16 .sum_lutc_input = "datac";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][6]~q ),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cycloneive_lcell_comb \mem~17 (
	.dataa(\mem[1][21]~q ),
	.datab(av_readdata_pre_21),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~17_combout ),
	.cout());
defparam \mem~17 .lut_mask = 16'hAACC;
defparam \mem~17 .sum_lutc_input = "datac";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][21]~q ),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cycloneive_lcell_comb \mem~18 (
	.dataa(\mem[1][30]~q ),
	.datab(av_readdata_pre_30),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~18_combout ),
	.cout());
defparam \mem~18 .lut_mask = 16'hAACC;
defparam \mem~18 .sum_lutc_input = "datac";

dffeas \mem[0][30] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][30]~q ),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[1][29] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

cycloneive_lcell_comb \mem~19 (
	.dataa(\mem[1][29]~q ),
	.datab(av_readdata_pre_29),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~19_combout ),
	.cout());
defparam \mem~19 .lut_mask = 16'hAACC;
defparam \mem~19 .sum_lutc_input = "datac";

dffeas \mem[0][29] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][29]~q ),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[1][28] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

cycloneive_lcell_comb \mem~20 (
	.dataa(\mem[1][28]~q ),
	.datab(av_readdata_pre_28),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~20_combout ),
	.cout());
defparam \mem~20 .lut_mask = 16'hAACC;
defparam \mem~20 .sum_lutc_input = "datac";

dffeas \mem[0][28] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][28]~q ),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[1][27] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

cycloneive_lcell_comb \mem~21 (
	.dataa(\mem[1][27]~q ),
	.datab(av_readdata_pre_27),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~21_combout ),
	.cout());
defparam \mem~21 .lut_mask = 16'hAACC;
defparam \mem~21 .sum_lutc_input = "datac";

dffeas \mem[0][27] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][27]~q ),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[1][26] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

cycloneive_lcell_comb \mem~22 (
	.dataa(\mem[1][26]~q ),
	.datab(av_readdata_pre_26),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~22_combout ),
	.cout());
defparam \mem~22 .lut_mask = 16'hAACC;
defparam \mem~22 .sum_lutc_input = "datac";

dffeas \mem[0][26] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][26]~q ),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[1][25] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

cycloneive_lcell_comb \mem~23 (
	.dataa(\mem[1][25]~q ),
	.datab(av_readdata_pre_25),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~23_combout ),
	.cout());
defparam \mem~23 .lut_mask = 16'hAACC;
defparam \mem~23 .sum_lutc_input = "datac";

dffeas \mem[0][25] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][25]~q ),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[1][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

cycloneive_lcell_comb \mem~24 (
	.dataa(\mem[1][24]~q ),
	.datab(av_readdata_pre_24),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~24_combout ),
	.cout());
defparam \mem~24 .lut_mask = 16'hAACC;
defparam \mem~24 .sum_lutc_input = "datac";

dffeas \mem[0][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][24]~q ),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[1][23] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

cycloneive_lcell_comb \mem~25 (
	.dataa(\mem[1][23]~q ),
	.datab(av_readdata_pre_23),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~25_combout ),
	.cout());
defparam \mem~25 .lut_mask = 16'hAACC;
defparam \mem~25 .sum_lutc_input = "datac";

dffeas \mem[0][23] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][23]~q ),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cycloneive_lcell_comb \mem~26 (
	.dataa(\mem[1][22]~q ),
	.datab(av_readdata_pre_22),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~26_combout ),
	.cout());
defparam \mem~26 .lut_mask = 16'hAACC;
defparam \mem~26 .sum_lutc_input = "datac";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][22]~q ),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cycloneive_lcell_comb \mem~27 (
	.dataa(\mem[1][20]~q ),
	.datab(av_readdata_pre_20),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~27_combout ),
	.cout());
defparam \mem~27 .lut_mask = 16'hAACC;
defparam \mem~27 .sum_lutc_input = "datac";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][20]~q ),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cycloneive_lcell_comb \mem~28 (
	.dataa(\mem[1][19]~q ),
	.datab(av_readdata_pre_19),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~28_combout ),
	.cout());
defparam \mem~28 .lut_mask = 16'hAACC;
defparam \mem~28 .sum_lutc_input = "datac";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][19]~q ),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cycloneive_lcell_comb \mem~29 (
	.dataa(\mem[1][18]~q ),
	.datab(av_readdata_pre_18),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~29_combout ),
	.cout());
defparam \mem~29 .lut_mask = 16'hAACC;
defparam \mem~29 .sum_lutc_input = "datac";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][18]~q ),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cycloneive_lcell_comb \mem~30 (
	.dataa(\mem[1][17]~q ),
	.datab(av_readdata_pre_17),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~30_combout ),
	.cout());
defparam \mem~30 .lut_mask = 16'hAACC;
defparam \mem~30 .sum_lutc_input = "datac";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][17]~q ),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[1][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

cycloneive_lcell_comb \mem~31 (
	.dataa(\mem[1][31]~q ),
	.datab(av_readdata_pre_31),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~31_combout ),
	.cout());
defparam \mem~31 .lut_mask = 16'hAACC;
defparam \mem~31 .sum_lutc_input = "datac";

dffeas \mem[0][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~4_combout ),
	.q(\mem[0][31]~q ),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

endmodule

module niosII_altera_avalon_sc_fifo_3 (
	clk,
	reset,
	saved_grant_1,
	mem_used_1,
	last_cycle,
	src_data_66,
	mem_used_0,
	mem_105_0,
	rp_valid,
	mem_84_0,
	mem_66_0,
	WideOr0,
	sink_ready,
	nonposted_write_endofpacket,
	uav_waitrequest,
	out_data_buffer_84,
	WideOr1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	saved_grant_1;
output 	mem_used_1;
input 	last_cycle;
input 	src_data_66;
output 	mem_used_0;
output 	mem_105_0;
input 	rp_valid;
output 	mem_84_0;
output 	mem_66_0;
input 	WideOr0;
input 	sink_ready;
input 	nonposted_write_endofpacket;
input 	uav_waitrequest;
input 	out_data_buffer_84;
input 	WideOr1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem_used[1]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~5_combout ;
wire \mem[1][105]~q ;
wire \mem~0_combout ;
wire \mem[1][84]~q ;
wire \mem~1_combout ;
wire \mem[1][66]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~2_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][84] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~2_combout ),
	.q(mem_84_0),
	.prn(vcc));
defparam \mem[0][84] .is_wysiwyg = "true";
defparam \mem[0][84] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~2_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(mem_used_0),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hAFFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~1 (
	.dataa(nonposted_write_endofpacket),
	.datab(WideOr1),
	.datac(src_data_66),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[0]~1_combout ),
	.cout());
defparam \mem_used[0]~1 .lut_mask = 16'hFEFE;
defparam \mem_used[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(mem_used_0),
	.datab(WideOr0),
	.datac(rp_valid),
	.datad(mem_105_0),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hFF7F;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~3 (
	.dataa(\mem_used[1]~0_combout ),
	.datab(\mem_used[0]~1_combout ),
	.datac(\mem_used[1]~2_combout ),
	.datad(uav_waitrequest),
	.cin(gnd),
	.combout(\mem_used[1]~3_combout ),
	.cout());
defparam \mem_used[1]~3 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(mem_used_0),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~5 (
	.dataa(\mem_used[0]~4_combout ),
	.datab(last_cycle),
	.datac(\mem_used[0]~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[0]~5_combout ),
	.cout());
defparam \mem_used[0]~5 .lut_mask = 16'hFEFE;
defparam \mem_used[0]~5 .sum_lutc_input = "datac";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][105]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

dffeas \mem[1][84] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][84]~q ),
	.prn(vcc));
defparam \mem[1][84] .is_wysiwyg = "true";
defparam \mem[1][84] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][84]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_84),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hFAFC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][66]~q ),
	.datab(src_data_66),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_4 (
	av_readdata_pre_22,
	av_readdata_pre_21,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_16,
	reset,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_105_0,
	mem_used_01,
	rp_valid,
	in_ready,
	av_readdata_pre_0,
	out_data_0,
	av_readdata_pre_1,
	out_data_1,
	av_readdata_pre_2,
	out_data_2,
	av_readdata_pre_3,
	out_data_3,
	av_readdata_pre_4,
	out_data_4,
	av_readdata_pre_5,
	out_data_5,
	av_readdata_pre_6,
	out_data_6,
	av_readdata_pre_7,
	out_data_7,
	out_data_22,
	out_data_21,
	out_data_20,
	out_data_19,
	out_data_18,
	out_data_17,
	out_data_16,
	av_readdata_pre_15,
	out_data_15,
	av_readdata_pre_14,
	out_data_14,
	av_readdata_pre_13,
	out_data_13,
	av_readdata_pre_12,
	out_data_12,
	av_readdata_pre_10,
	out_data_10,
	av_readdata_pre_9,
	out_data_9,
	av_readdata_pre_8,
	out_data_8,
	clk)/* synthesis synthesis_greybox=1 */;
input 	av_readdata_pre_22;
input 	av_readdata_pre_21;
input 	av_readdata_pre_20;
input 	av_readdata_pre_19;
input 	av_readdata_pre_18;
input 	av_readdata_pre_17;
input 	av_readdata_pre_16;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_105_0;
input 	mem_used_01;
input 	rp_valid;
input 	in_ready;
input 	av_readdata_pre_0;
output 	out_data_0;
input 	av_readdata_pre_1;
output 	out_data_1;
input 	av_readdata_pre_2;
output 	out_data_2;
input 	av_readdata_pre_3;
output 	out_data_3;
input 	av_readdata_pre_4;
output 	out_data_4;
input 	av_readdata_pre_5;
output 	out_data_5;
input 	av_readdata_pre_6;
output 	out_data_6;
input 	av_readdata_pre_7;
output 	out_data_7;
output 	out_data_22;
output 	out_data_21;
output 	out_data_20;
output 	out_data_19;
output 	out_data_18;
output 	out_data_17;
output 	out_data_16;
input 	av_readdata_pre_15;
output 	out_data_15;
input 	av_readdata_pre_14;
output 	out_data_14;
input 	av_readdata_pre_13;
output 	out_data_13;
input 	av_readdata_pre_12;
output 	out_data_12;
input 	av_readdata_pre_10;
output 	out_data_10;
input 	av_readdata_pre_9;
output 	out_data_9;
input 	av_readdata_pre_8;
output 	out_data_8;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[0][0]~q ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[0][1]~q ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[0][2]~q ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[0][3]~q ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[0][4]~q ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[0][5]~q ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[0][6]~q ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[0][7]~q ;
wire \mem[1][22]~q ;
wire \mem~8_combout ;
wire \mem[0][22]~q ;
wire \mem[1][21]~q ;
wire \mem~9_combout ;
wire \mem[0][21]~q ;
wire \mem[1][20]~q ;
wire \mem~10_combout ;
wire \mem[0][20]~q ;
wire \mem[1][19]~q ;
wire \mem~11_combout ;
wire \mem[0][19]~q ;
wire \mem[1][18]~q ;
wire \mem~12_combout ;
wire \mem[0][18]~q ;
wire \mem[1][17]~q ;
wire \mem~13_combout ;
wire \mem[0][17]~q ;
wire \mem[1][16]~q ;
wire \mem~14_combout ;
wire \mem[0][16]~q ;
wire \mem[1][15]~q ;
wire \mem~15_combout ;
wire \mem[0][15]~q ;
wire \mem[1][14]~q ;
wire \mem~16_combout ;
wire \mem[0][14]~q ;
wire \mem[1][13]~q ;
wire \mem~17_combout ;
wire \mem[0][13]~q ;
wire \mem[1][12]~q ;
wire \mem~18_combout ;
wire \mem[0][12]~q ;
wire \mem[1][10]~q ;
wire \mem~19_combout ;
wire \mem[0][10]~q ;
wire \mem[1][9]~q ;
wire \mem~20_combout ;
wire \mem[0][9]~q ;
wire \mem[1][8]~q ;
wire \mem~21_combout ;
wire \mem[0][8]~q ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \out_data[0]~0 (
	.dataa(\mem[0][0]~q ),
	.datab(av_readdata_pre_0),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_0),
	.cout());
defparam \out_data[0]~0 .lut_mask = 16'hEFFE;
defparam \out_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[1]~1 (
	.dataa(\mem[0][1]~q ),
	.datab(av_readdata_pre_1),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_1),
	.cout());
defparam \out_data[1]~1 .lut_mask = 16'hEFFE;
defparam \out_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[2]~2 (
	.dataa(\mem[0][2]~q ),
	.datab(av_readdata_pre_2),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_2),
	.cout());
defparam \out_data[2]~2 .lut_mask = 16'hEFFE;
defparam \out_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[3]~3 (
	.dataa(\mem[0][3]~q ),
	.datab(av_readdata_pre_3),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_3),
	.cout());
defparam \out_data[3]~3 .lut_mask = 16'hEFFE;
defparam \out_data[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[4]~4 (
	.dataa(\mem[0][4]~q ),
	.datab(av_readdata_pre_4),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_4),
	.cout());
defparam \out_data[4]~4 .lut_mask = 16'hEFFE;
defparam \out_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[5]~5 (
	.dataa(\mem[0][5]~q ),
	.datab(av_readdata_pre_5),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_5),
	.cout());
defparam \out_data[5]~5 .lut_mask = 16'hEFFE;
defparam \out_data[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[6]~6 (
	.dataa(\mem[0][6]~q ),
	.datab(av_readdata_pre_6),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_6),
	.cout());
defparam \out_data[6]~6 .lut_mask = 16'hEFFE;
defparam \out_data[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[7]~7 (
	.dataa(\mem[0][7]~q ),
	.datab(av_readdata_pre_7),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_7),
	.cout());
defparam \out_data[7]~7 .lut_mask = 16'hEFFE;
defparam \out_data[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[22]~8 (
	.dataa(\mem[0][22]~q ),
	.datab(av_readdata_pre_22),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_22),
	.cout());
defparam \out_data[22]~8 .lut_mask = 16'hEFFE;
defparam \out_data[22]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[21]~9 (
	.dataa(\mem[0][21]~q ),
	.datab(av_readdata_pre_21),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_21),
	.cout());
defparam \out_data[21]~9 .lut_mask = 16'hEFFE;
defparam \out_data[21]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[20]~10 (
	.dataa(\mem[0][20]~q ),
	.datab(av_readdata_pre_20),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_20),
	.cout());
defparam \out_data[20]~10 .lut_mask = 16'hEFFE;
defparam \out_data[20]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[19]~11 (
	.dataa(\mem[0][19]~q ),
	.datab(av_readdata_pre_19),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_19),
	.cout());
defparam \out_data[19]~11 .lut_mask = 16'hEFFE;
defparam \out_data[19]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[18]~12 (
	.dataa(\mem[0][18]~q ),
	.datab(av_readdata_pre_18),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_18),
	.cout());
defparam \out_data[18]~12 .lut_mask = 16'hEFFE;
defparam \out_data[18]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[17]~13 (
	.dataa(\mem[0][17]~q ),
	.datab(av_readdata_pre_17),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_17),
	.cout());
defparam \out_data[17]~13 .lut_mask = 16'hEFFE;
defparam \out_data[17]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[16]~14 (
	.dataa(\mem[0][16]~q ),
	.datab(av_readdata_pre_16),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_16),
	.cout());
defparam \out_data[16]~14 .lut_mask = 16'hEFFE;
defparam \out_data[16]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[15]~15 (
	.dataa(\mem[0][15]~q ),
	.datab(av_readdata_pre_15),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_15),
	.cout());
defparam \out_data[15]~15 .lut_mask = 16'hEFFE;
defparam \out_data[15]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[14]~16 (
	.dataa(\mem[0][14]~q ),
	.datab(av_readdata_pre_14),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_14),
	.cout());
defparam \out_data[14]~16 .lut_mask = 16'hEFFE;
defparam \out_data[14]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[13]~17 (
	.dataa(\mem[0][13]~q ),
	.datab(av_readdata_pre_13),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_13),
	.cout());
defparam \out_data[13]~17 .lut_mask = 16'hEFFE;
defparam \out_data[13]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[12]~18 (
	.dataa(\mem[0][12]~q ),
	.datab(av_readdata_pre_12),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_12),
	.cout());
defparam \out_data[12]~18 .lut_mask = 16'hEFFE;
defparam \out_data[12]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[10]~19 (
	.dataa(\mem[0][10]~q ),
	.datab(av_readdata_pre_10),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_10),
	.cout());
defparam \out_data[10]~19 .lut_mask = 16'hEFFE;
defparam \out_data[10]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[9]~20 (
	.dataa(\mem[0][9]~q ),
	.datab(av_readdata_pre_9),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_9),
	.cout());
defparam \out_data[9]~20 .lut_mask = 16'hEFFE;
defparam \out_data[9]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[8]~21 (
	.dataa(\mem[0][8]~q ),
	.datab(av_readdata_pre_8),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(out_data_8),
	.cout());
defparam \out_data[8]~21 .lut_mask = 16'hEFFE;
defparam \out_data[8]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(mem_105_0),
	.datab(mem_used_01),
	.datac(rp_valid),
	.datad(in_ready),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h7FFF;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[1]~q ),
	.datab(read_latency_shift_reg_0),
	.datac(mem_used_0),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~0 (
	.dataa(\mem_used[1]~q ),
	.datab(mem_used_0),
	.datac(read_latency_shift_reg_0),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~0_combout ),
	.cout());
defparam \mem_used[0]~0 .lut_mask = 16'hFDFE;
defparam \mem_used[0]~0 .sum_lutc_input = "datac";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][0]~q ),
	.datab(av_readdata_pre_0),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hAAFF;
defparam \always0~0 .sum_lutc_input = "datac";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][0]~q ),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][1]~q ),
	.datab(av_readdata_pre_1),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][1]~q ),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][2]~q ),
	.datab(av_readdata_pre_2),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][2]~q ),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][3]~q ),
	.datab(av_readdata_pre_3),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hAACC;
defparam \mem~3 .sum_lutc_input = "datac";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][3]~q ),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[1][4]~q ),
	.datab(av_readdata_pre_4),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hAACC;
defparam \mem~4 .sum_lutc_input = "datac";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][4]~q ),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cycloneive_lcell_comb \mem~5 (
	.dataa(\mem[1][5]~q ),
	.datab(av_readdata_pre_5),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~5_combout ),
	.cout());
defparam \mem~5 .lut_mask = 16'hAACC;
defparam \mem~5 .sum_lutc_input = "datac";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][5]~q ),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cycloneive_lcell_comb \mem~6 (
	.dataa(\mem[1][6]~q ),
	.datab(av_readdata_pre_6),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~6_combout ),
	.cout());
defparam \mem~6 .lut_mask = 16'hAACC;
defparam \mem~6 .sum_lutc_input = "datac";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][6]~q ),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cycloneive_lcell_comb \mem~7 (
	.dataa(\mem[1][7]~q ),
	.datab(av_readdata_pre_7),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~7_combout ),
	.cout());
defparam \mem~7 .lut_mask = 16'hAACC;
defparam \mem~7 .sum_lutc_input = "datac";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][7]~q ),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cycloneive_lcell_comb \mem~8 (
	.dataa(\mem[1][22]~q ),
	.datab(av_readdata_pre_22),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~8_combout ),
	.cout());
defparam \mem~8 .lut_mask = 16'hAACC;
defparam \mem~8 .sum_lutc_input = "datac";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][22]~q ),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cycloneive_lcell_comb \mem~9 (
	.dataa(\mem[1][21]~q ),
	.datab(av_readdata_pre_21),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~9_combout ),
	.cout());
defparam \mem~9 .lut_mask = 16'hAACC;
defparam \mem~9 .sum_lutc_input = "datac";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][21]~q ),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cycloneive_lcell_comb \mem~10 (
	.dataa(\mem[1][20]~q ),
	.datab(av_readdata_pre_20),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~10_combout ),
	.cout());
defparam \mem~10 .lut_mask = 16'hAACC;
defparam \mem~10 .sum_lutc_input = "datac";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][20]~q ),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cycloneive_lcell_comb \mem~11 (
	.dataa(\mem[1][19]~q ),
	.datab(av_readdata_pre_19),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~11_combout ),
	.cout());
defparam \mem~11 .lut_mask = 16'hAACC;
defparam \mem~11 .sum_lutc_input = "datac";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][19]~q ),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cycloneive_lcell_comb \mem~12 (
	.dataa(\mem[1][18]~q ),
	.datab(av_readdata_pre_18),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~12_combout ),
	.cout());
defparam \mem~12 .lut_mask = 16'hAACC;
defparam \mem~12 .sum_lutc_input = "datac";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][18]~q ),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cycloneive_lcell_comb \mem~13 (
	.dataa(\mem[1][17]~q ),
	.datab(av_readdata_pre_17),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~13_combout ),
	.cout());
defparam \mem~13 .lut_mask = 16'hAACC;
defparam \mem~13 .sum_lutc_input = "datac";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][17]~q ),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cycloneive_lcell_comb \mem~14 (
	.dataa(\mem[1][16]~q ),
	.datab(av_readdata_pre_16),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~14_combout ),
	.cout());
defparam \mem~14 .lut_mask = 16'hAACC;
defparam \mem~14 .sum_lutc_input = "datac";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][16]~q ),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cycloneive_lcell_comb \mem~15 (
	.dataa(\mem[1][15]~q ),
	.datab(av_readdata_pre_15),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~15_combout ),
	.cout());
defparam \mem~15 .lut_mask = 16'hAACC;
defparam \mem~15 .sum_lutc_input = "datac";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][15]~q ),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cycloneive_lcell_comb \mem~16 (
	.dataa(\mem[1][14]~q ),
	.datab(av_readdata_pre_14),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~16_combout ),
	.cout());
defparam \mem~16 .lut_mask = 16'hAACC;
defparam \mem~16 .sum_lutc_input = "datac";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][14]~q ),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cycloneive_lcell_comb \mem~17 (
	.dataa(\mem[1][13]~q ),
	.datab(av_readdata_pre_13),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~17_combout ),
	.cout());
defparam \mem~17 .lut_mask = 16'hAACC;
defparam \mem~17 .sum_lutc_input = "datac";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][13]~q ),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cycloneive_lcell_comb \mem~18 (
	.dataa(\mem[1][12]~q ),
	.datab(av_readdata_pre_12),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~18_combout ),
	.cout());
defparam \mem~18 .lut_mask = 16'hAACC;
defparam \mem~18 .sum_lutc_input = "datac";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][12]~q ),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cycloneive_lcell_comb \mem~19 (
	.dataa(\mem[1][10]~q ),
	.datab(av_readdata_pre_10),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~19_combout ),
	.cout());
defparam \mem~19 .lut_mask = 16'hAACC;
defparam \mem~19 .sum_lutc_input = "datac";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][10]~q ),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cycloneive_lcell_comb \mem~20 (
	.dataa(\mem[1][9]~q ),
	.datab(av_readdata_pre_9),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~20_combout ),
	.cout());
defparam \mem~20 .lut_mask = 16'hAACC;
defparam \mem~20 .sum_lutc_input = "datac";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][9]~q ),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cycloneive_lcell_comb \mem~21 (
	.dataa(\mem[1][8]~q ),
	.datab(av_readdata_pre_8),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~21_combout ),
	.cout());
defparam \mem~21 .lut_mask = 16'hAACC;
defparam \mem~21 .sum_lutc_input = "datac";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][8]~q ),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

endmodule

module niosII_altera_avalon_sc_fifo_5 (
	reset,
	in_data_toggle,
	out_data_toggle_flopped,
	dreg_0,
	mem_used_1,
	out_data_buffer_66,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_105_0,
	mem_used_01,
	dreg_01,
	out_data_buffer_65,
	read_latency_shift_reg,
	out_data_buffer_105,
	out_data_buffer_64,
	in_ready,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	in_data_toggle;
input 	out_data_toggle_flopped;
input 	dreg_0;
output 	mem_used_1;
input 	out_data_buffer_66;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
output 	mem_105_0;
output 	mem_used_01;
input 	dreg_01;
input 	out_data_buffer_65;
input 	read_latency_shift_reg;
input 	out_data_buffer_105;
input 	out_data_buffer_64;
input 	in_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem~0_combout ;
wire \write~0_combout ;
wire \read~4_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[0][105]~1_combout ;
wire \mem~2_combout ;
wire \mem[1][105]~q ;
wire \mem~3_combout ;
wire \mem[0][105]~4_combout ;
wire \mem_used[0]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem[0][105]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_01),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(out_data_buffer_65),
	.datab(out_data_buffer_105),
	.datac(gnd),
	.datad(out_data_buffer_64),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hEEFF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~0 (
	.dataa(read_latency_shift_reg),
	.datab(out_data_buffer_66),
	.datac(\mem~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFEFE;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~4 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_used_0),
	.datac(mem_105_0),
	.datad(in_ready),
	.cin(gnd),
	.combout(\read~4_combout ),
	.cout());
defparam \read~4 .lut_mask = 16'hFEFF;
defparam \read~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(mem_used_1),
	.datab(mem_used_01),
	.datac(\write~0_combout ),
	.datad(\read~4_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hBEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][105]~1 (
	.dataa(mem_105_0),
	.datab(mem_used_01),
	.datac(in_data_toggle),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\mem[0][105]~1_combout ),
	.cout());
defparam \mem[0][105]~1 .lut_mask = 16'hEFFE;
defparam \mem[0][105]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~2 (
	.dataa(gnd),
	.datab(out_data_toggle_flopped),
	.datac(dreg_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'h3CFF;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(mem_used_1),
	.datab(\mem~2_combout ),
	.datac(\mem~0_combout ),
	.datad(\mem[1][105]~q ),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hFFFE;
defparam \mem~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][105]~4 (
	.dataa(\mem[0][105]~1_combout ),
	.datab(\mem~3_combout ),
	.datac(\read~4_combout ),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(\mem[0][105]~4_combout ),
	.cout());
defparam \mem[0][105]~4 .lut_mask = 16'hFEFF;
defparam \mem[0][105]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~1 (
	.dataa(\write~0_combout ),
	.datab(mem_used_01),
	.datac(mem_used_1),
	.datad(\read~4_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~1_combout ),
	.cout());
defparam \mem_used[0]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_6 (
	clk,
	reset,
	uav_read,
	hold_waitrequest,
	Equal6,
	src_channel_12,
	read_latency_shift_reg_0,
	mem_used_1,
	read_latency_shift_reg)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	uav_read;
input 	hold_waitrequest;
input 	Equal6;
input 	src_channel_12;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	read_latency_shift_reg;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(hold_waitrequest),
	.datab(uav_read),
	.datac(Equal6),
	.datad(src_channel_12),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFFFE;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_7 (
	clk,
	W_alu_result_5,
	W_alu_result_4,
	reset,
	d_read,
	read_accepted,
	uav_read,
	hold_waitrequest,
	cp_valid,
	src_channel_12,
	read_latency_shift_reg_0,
	mem_used_1,
	write)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	reset;
input 	d_read;
input 	read_accepted;
input 	uav_read;
input 	hold_waitrequest;
input 	cp_valid;
input 	src_channel_12;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
output 	write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(W_alu_result_5),
	.datab(W_alu_result_4),
	.datac(src_channel_12),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(write),
	.cout());
defparam \write~0 .lut_mask = 16'hFEFF;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(uav_read),
	.datac(cp_valid),
	.datad(write),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(W_alu_result_5),
	.datab(hold_waitrequest),
	.datac(read_accepted),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hEFEF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(W_alu_result_4),
	.datab(src_channel_12),
	.datac(d_read),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFFFE;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~1_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_8 (
	clk,
	reset,
	uav_read,
	hold_waitrequest,
	Equal9,
	mem_used_1,
	Equal5,
	read_latency_shift_reg_0,
	read_latency_shift_reg)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	uav_read;
input 	hold_waitrequest;
input 	Equal9;
output 	mem_used_1;
input 	Equal5;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(hold_waitrequest),
	.datab(uav_read),
	.datac(Equal9),
	.datad(Equal5),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFFFE;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_9 (
	clk,
	W_alu_result_5,
	W_alu_result_4,
	reset,
	d_read,
	read_accepted,
	uav_read,
	hold_waitrequest,
	cp_valid,
	src_channel_12,
	read_latency_shift_reg_0,
	write,
	write1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	reset;
input 	d_read;
input 	read_accepted;
input 	uav_read;
input 	hold_waitrequest;
input 	cp_valid;
input 	src_channel_12;
input 	read_latency_shift_reg_0;
output 	write;
output 	write1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem_used[1]~q ;


cycloneive_lcell_comb \write~2 (
	.dataa(W_alu_result_5),
	.datab(src_channel_12),
	.datac(W_alu_result_4),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(write),
	.cout());
defparam \write~2 .lut_mask = 16'hEFFF;
defparam \write~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~3 (
	.dataa(d_read),
	.datab(read_accepted),
	.datac(hold_waitrequest),
	.datad(gnd),
	.cin(gnd),
	.combout(write1),
	.cout());
defparam \write~3 .lut_mask = 16'hFBFB;
defparam \write~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(\mem_used[1]~q ),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(uav_read),
	.datac(cp_valid),
	.datad(write),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(hold_waitrequest),
	.datab(uav_read),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(W_alu_result_5),
	.datab(src_channel_12),
	.datac(\mem_used[1]~0_combout ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(\mem_used[1]~q ),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

endmodule

module niosII_altera_avalon_sc_fifo_10 (
	clk,
	reset,
	read_latency_shift_reg_0,
	Equal12,
	mem_used_1,
	read_latency_shift_reg,
	read_latency_shift_reg1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	read_latency_shift_reg_0;
input 	Equal12;
output 	mem_used_1;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(read_latency_shift_reg1),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(Equal12),
	.datab(read_latency_shift_reg),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[1]~0_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_11 (
	clk,
	W_alu_result_3,
	reset,
	uav_read,
	hold_waitrequest,
	Equal9,
	Equal6,
	read_latency_shift_reg_0,
	mem_used_1,
	read_latency_shift_reg)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_3;
input 	reset;
input 	uav_read;
input 	hold_waitrequest;
input 	Equal9;
input 	Equal6;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	read_latency_shift_reg;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(hold_waitrequest),
	.datab(uav_read),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(W_alu_result_3),
	.datab(Equal9),
	.datac(Equal6),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFFFE;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_12 (
	clk,
	reset,
	out_valid1,
	mem_used_0,
	mem_87_0,
	out_payload_0,
	out_payload_1,
	out_payload_2,
	out_payload_3,
	out_payload_4,
	out_payload_11,
	out_payload_13,
	out_payload_12,
	out_payload_5,
	out_payload_14,
	out_payload_15,
	out_payload_10,
	out_payload_9,
	out_payload_8,
	out_payload_7,
	out_payload_6,
	za_valid,
	za_data_0,
	za_data_1,
	za_data_2,
	za_data_3,
	za_data_4,
	za_data_11,
	za_data_13,
	za_data_12,
	za_data_5,
	za_data_14,
	za_data_15,
	za_data_10,
	za_data_9,
	za_data_8,
	za_data_7,
	za_data_6)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
output 	out_valid1;
input 	mem_used_0;
input 	mem_87_0;
output 	out_payload_0;
output 	out_payload_1;
output 	out_payload_2;
output 	out_payload_3;
output 	out_payload_4;
output 	out_payload_11;
output 	out_payload_13;
output 	out_payload_12;
output 	out_payload_5;
output 	out_payload_14;
output 	out_payload_15;
output 	out_payload_10;
output 	out_payload_9;
output 	out_payload_8;
output 	out_payload_7;
output 	out_payload_6;
input 	za_valid;
input 	za_data_0;
input 	za_data_1;
input 	za_data_2;
input 	za_data_3;
input 	za_data_4;
input 	za_data_11;
input 	za_data_13;
input 	za_data_12;
input 	za_data_5;
input 	za_data_14;
input 	za_data_15;
input 	za_data_10;
input 	za_data_9;
input 	za_data_8;
input 	za_data_7;
input 	za_data_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \internal_out_ready~0_combout ;
wire \mem_rd_ptr[0]~1_combout ;
wire \rd_ptr[0]~q ;
wire \mem_rd_ptr[1]~0_combout ;
wire \rd_ptr[1]~q ;
wire \wr_ptr[0]~0_combout ;
wire \next_full~2_combout ;
wire \mem_rd_ptr[2]~2_combout ;
wire \rd_ptr[2]~q ;
wire \wr_ptr[2]~q ;
wire \Add0~1_combout ;
wire \next_full~3_combout ;
wire \next_full~4_combout ;
wire \full~q ;
wire \write~combout ;
wire \wr_ptr[0]~q ;
wire \Add0~0_combout ;
wire \wr_ptr[1]~q ;
wire \internal_out_valid~0_combout ;
wire \Equal0~0_combout ;
wire \internal_out_valid~2_combout ;
wire \next_empty~0_combout ;
wire \empty~q ;
wire \internal_out_valid~1_combout ;
wire \internal_out_valid~q ;
wire \mem~208_combout ;
wire \mem~80_q ;
wire \mem~209_combout ;
wire \mem~96_q ;
wire \mem~210_combout ;
wire \mem~64_q ;
wire \mem~128_combout ;
wire \mem~211_combout ;
wire \mem~112_q ;
wire \mem~129_combout ;
wire \mem~212_combout ;
wire \mem~32_q ;
wire \mem~213_combout ;
wire \mem~16_q ;
wire \mem~214_combout ;
wire \mem~0_q ;
wire \mem~130_combout ;
wire \mem~215_combout ;
wire \mem~48_q ;
wire \mem~131_combout ;
wire \mem~132_combout ;
wire \internal_out_payload[0]~q ;
wire \mem~81_q ;
wire \mem~97_q ;
wire \mem~65_q ;
wire \mem~133_combout ;
wire \mem~113_q ;
wire \mem~134_combout ;
wire \mem~33_q ;
wire \mem~17_q ;
wire \mem~1_q ;
wire \mem~135_combout ;
wire \mem~49_q ;
wire \mem~136_combout ;
wire \mem~137_combout ;
wire \internal_out_payload[1]~q ;
wire \mem~82_q ;
wire \mem~98_q ;
wire \mem~66_q ;
wire \mem~138_combout ;
wire \mem~114_q ;
wire \mem~139_combout ;
wire \mem~34_q ;
wire \mem~18_q ;
wire \mem~2_q ;
wire \mem~140_combout ;
wire \mem~50_q ;
wire \mem~141_combout ;
wire \mem~142_combout ;
wire \internal_out_payload[2]~q ;
wire \mem~83_q ;
wire \mem~99_q ;
wire \mem~67_q ;
wire \mem~143_combout ;
wire \mem~115_q ;
wire \mem~144_combout ;
wire \mem~35_q ;
wire \mem~19_q ;
wire \mem~3_q ;
wire \mem~145_combout ;
wire \mem~51_q ;
wire \mem~146_combout ;
wire \mem~147_combout ;
wire \internal_out_payload[3]~q ;
wire \mem~84_q ;
wire \mem~100_q ;
wire \mem~68_q ;
wire \mem~148_combout ;
wire \mem~116_q ;
wire \mem~149_combout ;
wire \mem~36_q ;
wire \mem~20_q ;
wire \mem~4_q ;
wire \mem~150_combout ;
wire \mem~52_q ;
wire \mem~151_combout ;
wire \mem~152_combout ;
wire \internal_out_payload[4]~q ;
wire \mem~91_q ;
wire \mem~107_q ;
wire \mem~75_q ;
wire \mem~153_combout ;
wire \mem~123_q ;
wire \mem~154_combout ;
wire \mem~43_q ;
wire \mem~27_q ;
wire \mem~11_q ;
wire \mem~155_combout ;
wire \mem~59_q ;
wire \mem~156_combout ;
wire \mem~157_combout ;
wire \internal_out_payload[11]~q ;
wire \mem~93_q ;
wire \mem~109_q ;
wire \mem~77_q ;
wire \mem~158_combout ;
wire \mem~125_q ;
wire \mem~159_combout ;
wire \mem~45_q ;
wire \mem~29_q ;
wire \mem~13_q ;
wire \mem~160_combout ;
wire \mem~61_q ;
wire \mem~161_combout ;
wire \mem~162_combout ;
wire \internal_out_payload[13]~q ;
wire \mem~92_q ;
wire \mem~108_q ;
wire \mem~76_q ;
wire \mem~163_combout ;
wire \mem~124_q ;
wire \mem~164_combout ;
wire \mem~44_q ;
wire \mem~28_q ;
wire \mem~12_q ;
wire \mem~165_combout ;
wire \mem~60_q ;
wire \mem~166_combout ;
wire \mem~167_combout ;
wire \internal_out_payload[12]~q ;
wire \mem~85_q ;
wire \mem~101_q ;
wire \mem~69_q ;
wire \mem~168_combout ;
wire \mem~117_q ;
wire \mem~169_combout ;
wire \mem~37_q ;
wire \mem~21_q ;
wire \mem~5_q ;
wire \mem~170_combout ;
wire \mem~53_q ;
wire \mem~171_combout ;
wire \mem~172_combout ;
wire \internal_out_payload[5]~q ;
wire \mem~94_q ;
wire \mem~110_q ;
wire \mem~78_q ;
wire \mem~173_combout ;
wire \mem~126_q ;
wire \mem~174_combout ;
wire \mem~46_q ;
wire \mem~30_q ;
wire \mem~14_q ;
wire \mem~175_combout ;
wire \mem~62_q ;
wire \mem~176_combout ;
wire \mem~177_combout ;
wire \internal_out_payload[14]~q ;
wire \mem~95_q ;
wire \mem~111_q ;
wire \mem~79_q ;
wire \mem~178_combout ;
wire \mem~127_q ;
wire \mem~179_combout ;
wire \mem~47_q ;
wire \mem~31_q ;
wire \mem~15_q ;
wire \mem~180_combout ;
wire \mem~63_q ;
wire \mem~181_combout ;
wire \mem~182_combout ;
wire \internal_out_payload[15]~q ;
wire \mem~90_q ;
wire \mem~106_q ;
wire \mem~74_q ;
wire \mem~183_combout ;
wire \mem~122_q ;
wire \mem~184_combout ;
wire \mem~42_q ;
wire \mem~26_q ;
wire \mem~10_q ;
wire \mem~185_combout ;
wire \mem~58_q ;
wire \mem~186_combout ;
wire \mem~187_combout ;
wire \internal_out_payload[10]~q ;
wire \mem~89_q ;
wire \mem~105_q ;
wire \mem~73_q ;
wire \mem~188_combout ;
wire \mem~121_q ;
wire \mem~189_combout ;
wire \mem~41_q ;
wire \mem~25_q ;
wire \mem~9_q ;
wire \mem~190_combout ;
wire \mem~57_q ;
wire \mem~191_combout ;
wire \mem~192_combout ;
wire \internal_out_payload[9]~q ;
wire \mem~88_q ;
wire \mem~104_q ;
wire \mem~72_q ;
wire \mem~193_combout ;
wire \mem~120_q ;
wire \mem~194_combout ;
wire \mem~40_q ;
wire \mem~24_q ;
wire \mem~8_q ;
wire \mem~195_combout ;
wire \mem~56_q ;
wire \mem~196_combout ;
wire \mem~197_combout ;
wire \internal_out_payload[8]~q ;
wire \mem~87_q ;
wire \mem~103_q ;
wire \mem~71_q ;
wire \mem~198_combout ;
wire \mem~119_q ;
wire \mem~199_combout ;
wire \mem~39_q ;
wire \mem~23_q ;
wire \mem~7_q ;
wire \mem~200_combout ;
wire \mem~55_q ;
wire \mem~201_combout ;
wire \mem~202_combout ;
wire \internal_out_payload[7]~q ;
wire \mem~86_q ;
wire \mem~102_q ;
wire \mem~70_q ;
wire \mem~203_combout ;
wire \mem~118_q ;
wire \mem~204_combout ;
wire \mem~38_q ;
wire \mem~22_q ;
wire \mem~6_q ;
wire \mem~205_combout ;
wire \mem~54_q ;
wire \mem~206_combout ;
wire \mem~207_combout ;
wire \internal_out_payload[6]~q ;


dffeas out_valid(
	.clk(clk),
	.d(\internal_out_valid~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_payload[0] (
	.clk(clk),
	.d(\internal_out_payload[0]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_0),
	.prn(vcc));
defparam \out_payload[0] .is_wysiwyg = "true";
defparam \out_payload[0] .power_up = "low";

dffeas \out_payload[1] (
	.clk(clk),
	.d(\internal_out_payload[1]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_1),
	.prn(vcc));
defparam \out_payload[1] .is_wysiwyg = "true";
defparam \out_payload[1] .power_up = "low";

dffeas \out_payload[2] (
	.clk(clk),
	.d(\internal_out_payload[2]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_2),
	.prn(vcc));
defparam \out_payload[2] .is_wysiwyg = "true";
defparam \out_payload[2] .power_up = "low";

dffeas \out_payload[3] (
	.clk(clk),
	.d(\internal_out_payload[3]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_3),
	.prn(vcc));
defparam \out_payload[3] .is_wysiwyg = "true";
defparam \out_payload[3] .power_up = "low";

dffeas \out_payload[4] (
	.clk(clk),
	.d(\internal_out_payload[4]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_4),
	.prn(vcc));
defparam \out_payload[4] .is_wysiwyg = "true";
defparam \out_payload[4] .power_up = "low";

dffeas \out_payload[11] (
	.clk(clk),
	.d(\internal_out_payload[11]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_11),
	.prn(vcc));
defparam \out_payload[11] .is_wysiwyg = "true";
defparam \out_payload[11] .power_up = "low";

dffeas \out_payload[13] (
	.clk(clk),
	.d(\internal_out_payload[13]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_13),
	.prn(vcc));
defparam \out_payload[13] .is_wysiwyg = "true";
defparam \out_payload[13] .power_up = "low";

dffeas \out_payload[12] (
	.clk(clk),
	.d(\internal_out_payload[12]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_12),
	.prn(vcc));
defparam \out_payload[12] .is_wysiwyg = "true";
defparam \out_payload[12] .power_up = "low";

dffeas \out_payload[5] (
	.clk(clk),
	.d(\internal_out_payload[5]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_5),
	.prn(vcc));
defparam \out_payload[5] .is_wysiwyg = "true";
defparam \out_payload[5] .power_up = "low";

dffeas \out_payload[14] (
	.clk(clk),
	.d(\internal_out_payload[14]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_14),
	.prn(vcc));
defparam \out_payload[14] .is_wysiwyg = "true";
defparam \out_payload[14] .power_up = "low";

dffeas \out_payload[15] (
	.clk(clk),
	.d(\internal_out_payload[15]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_15),
	.prn(vcc));
defparam \out_payload[15] .is_wysiwyg = "true";
defparam \out_payload[15] .power_up = "low";

dffeas \out_payload[10] (
	.clk(clk),
	.d(\internal_out_payload[10]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_10),
	.prn(vcc));
defparam \out_payload[10] .is_wysiwyg = "true";
defparam \out_payload[10] .power_up = "low";

dffeas \out_payload[9] (
	.clk(clk),
	.d(\internal_out_payload[9]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_9),
	.prn(vcc));
defparam \out_payload[9] .is_wysiwyg = "true";
defparam \out_payload[9] .power_up = "low";

dffeas \out_payload[8] (
	.clk(clk),
	.d(\internal_out_payload[8]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_8),
	.prn(vcc));
defparam \out_payload[8] .is_wysiwyg = "true";
defparam \out_payload[8] .power_up = "low";

dffeas \out_payload[7] (
	.clk(clk),
	.d(\internal_out_payload[7]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_7),
	.prn(vcc));
defparam \out_payload[7] .is_wysiwyg = "true";
defparam \out_payload[7] .power_up = "low";

dffeas \out_payload[6] (
	.clk(clk),
	.d(\internal_out_payload[6]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_6),
	.prn(vcc));
defparam \out_payload[6] .is_wysiwyg = "true";
defparam \out_payload[6] .power_up = "low";

cycloneive_lcell_comb \read~0 (
	.dataa(\internal_out_valid~q ),
	.datab(mem_used_0),
	.datac(mem_87_0),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hBFFF;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_out_ready~0 (
	.dataa(gnd),
	.datab(mem_used_0),
	.datac(mem_87_0),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\internal_out_ready~0_combout ),
	.cout());
defparam \internal_out_ready~0 .lut_mask = 16'h3FFF;
defparam \internal_out_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[0]~1 (
	.dataa(gnd),
	.datab(\rd_ptr[0]~q ),
	.datac(\internal_out_valid~q ),
	.datad(\internal_out_ready~0_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[0]~1_combout ),
	.cout());
defparam \mem_rd_ptr[0]~1 .lut_mask = 16'hC33C;
defparam \mem_rd_ptr[0]~1 .sum_lutc_input = "datac";

dffeas \rd_ptr[0] (
	.clk(clk),
	.d(\mem_rd_ptr[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[0]~q ),
	.prn(vcc));
defparam \rd_ptr[0] .is_wysiwyg = "true";
defparam \rd_ptr[0] .power_up = "low";

cycloneive_lcell_comb \mem_rd_ptr[1]~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\internal_out_valid~q ),
	.datac(\internal_out_ready~0_combout ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[1]~0_combout ),
	.cout());
defparam \mem_rd_ptr[1]~0 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[1]~0 .sum_lutc_input = "datac";

dffeas \rd_ptr[1] (
	.clk(clk),
	.d(\mem_rd_ptr[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[1]~q ),
	.prn(vcc));
defparam \rd_ptr[1] .is_wysiwyg = "true";
defparam \rd_ptr[1] .power_up = "low";

cycloneive_lcell_comb \wr_ptr[0]~0 (
	.dataa(\wr_ptr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_ptr[0]~0_combout ),
	.cout());
defparam \wr_ptr[0]~0 .lut_mask = 16'h5555;
defparam \wr_ptr[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~2 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\rd_ptr[0]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\next_full~2_combout ),
	.cout());
defparam \next_full~2 .lut_mask = 16'h6996;
defparam \next_full~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[2]~2 (
	.dataa(\rd_ptr[2]~q ),
	.datab(\read~0_combout ),
	.datac(\rd_ptr[1]~q ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[2]~2_combout ),
	.cout());
defparam \mem_rd_ptr[2]~2 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[2]~2 .sum_lutc_input = "datac";

dffeas \rd_ptr[2] (
	.clk(clk),
	.d(\mem_rd_ptr[2]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[2]~q ),
	.prn(vcc));
defparam \rd_ptr[2] .is_wysiwyg = "true";
defparam \rd_ptr[2] .power_up = "low";

dffeas \wr_ptr[2] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[2]~q ),
	.prn(vcc));
defparam \wr_ptr[2] .is_wysiwyg = "true";
defparam \wr_ptr[2] .power_up = "low";

cycloneive_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'hC33C;
defparam \Add0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~3 (
	.dataa(\next_full~2_combout ),
	.datab(\rd_ptr[2]~q ),
	.datac(\Add0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_full~3_combout ),
	.cout());
defparam \next_full~3 .lut_mask = 16'hBEBE;
defparam \next_full~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~4 (
	.dataa(za_valid),
	.datab(\full~q ),
	.datac(\next_full~3_combout ),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\next_full~4_combout ),
	.cout());
defparam \next_full~4 .lut_mask = 16'hFEFF;
defparam \next_full~4 .sum_lutc_input = "datac";

dffeas full(
	.clk(clk),
	.d(\next_full~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\full~q ),
	.prn(vcc));
defparam full.is_wysiwyg = "true";
defparam full.power_up = "low";

cycloneive_lcell_comb write(
	.dataa(za_valid),
	.datab(gnd),
	.datac(gnd),
	.datad(\full~q ),
	.cin(gnd),
	.combout(\write~combout ),
	.cout());
defparam write.lut_mask = 16'hAAFF;
defparam write.sum_lutc_input = "datac";

dffeas \wr_ptr[0] (
	.clk(clk),
	.d(\wr_ptr[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[0]~q ),
	.prn(vcc));
defparam \wr_ptr[0] .is_wysiwyg = "true";
defparam \wr_ptr[0] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h0FF0;
defparam \Add0~0 .sum_lutc_input = "datac";

dffeas \wr_ptr[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[1]~q ),
	.prn(vcc));
defparam \wr_ptr[1] .is_wysiwyg = "true";
defparam \wr_ptr[1] .power_up = "low";

cycloneive_lcell_comb \internal_out_valid~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\internal_out_valid~0_combout ),
	.cout());
defparam \internal_out_valid~0 .lut_mask = 16'h6996;
defparam \internal_out_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\rd_ptr[0]~q ),
	.datac(\wr_ptr[2]~q ),
	.datad(\rd_ptr[2]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_out_valid~2 (
	.dataa(\internal_out_valid~q ),
	.datab(\internal_out_ready~0_combout ),
	.datac(\internal_out_valid~0_combout ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\internal_out_valid~2_combout ),
	.cout());
defparam \internal_out_valid~2 .lut_mask = 16'hFEFF;
defparam \internal_out_valid~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_empty~0 (
	.dataa(\read~0_combout ),
	.datab(\internal_out_valid~2_combout ),
	.datac(\empty~q ),
	.datad(\write~combout ),
	.cin(gnd),
	.combout(\next_empty~0_combout ),
	.cout());
defparam \next_empty~0 .lut_mask = 16'hFFF7;
defparam \next_empty~0 .sum_lutc_input = "datac";

dffeas empty(
	.clk(clk),
	.d(\next_empty~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty~q ),
	.prn(vcc));
defparam empty.is_wysiwyg = "true";
defparam empty.power_up = "low";

cycloneive_lcell_comb \internal_out_valid~1 (
	.dataa(\read~0_combout ),
	.datab(\internal_out_valid~0_combout ),
	.datac(\Equal0~0_combout ),
	.datad(\empty~q ),
	.cin(gnd),
	.combout(\internal_out_valid~1_combout ),
	.cout());
defparam \internal_out_valid~1 .lut_mask = 16'hFFF7;
defparam \internal_out_valid~1 .sum_lutc_input = "datac";

dffeas internal_out_valid(
	.clk(clk),
	.d(\internal_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_valid~q ),
	.prn(vcc));
defparam internal_out_valid.is_wysiwyg = "true";
defparam internal_out_valid.power_up = "low";

cycloneive_lcell_comb \mem~208 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\wr_ptr[0]~q ),
	.datac(\write~combout ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~208_combout ),
	.cout());
defparam \mem~208 .lut_mask = 16'hFEFF;
defparam \mem~208 .sum_lutc_input = "datac";

dffeas \mem~80 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~80_q ),
	.prn(vcc));
defparam \mem~80 .is_wysiwyg = "true";
defparam \mem~80 .power_up = "low";

cycloneive_lcell_comb \mem~209 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\write~combout ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem~209_combout ),
	.cout());
defparam \mem~209 .lut_mask = 16'hFEFF;
defparam \mem~209 .sum_lutc_input = "datac";

dffeas \mem~96 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~96_q ),
	.prn(vcc));
defparam \mem~96 .is_wysiwyg = "true";
defparam \mem~96 .power_up = "low";

cycloneive_lcell_comb \mem~210 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\write~combout ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~210_combout ),
	.cout());
defparam \mem~210 .lut_mask = 16'hEFFF;
defparam \mem~210 .sum_lutc_input = "datac";

dffeas \mem~64 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~64_q ),
	.prn(vcc));
defparam \mem~64 .is_wysiwyg = "true";
defparam \mem~64 .power_up = "low";

cycloneive_lcell_comb \mem~128 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~96_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~64_q ),
	.cin(gnd),
	.combout(\mem~128_combout ),
	.cout());
defparam \mem~128 .lut_mask = 16'hFFDE;
defparam \mem~128 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~211 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\wr_ptr[0]~q ),
	.datac(\wr_ptr[1]~q ),
	.datad(\write~combout ),
	.cin(gnd),
	.combout(\mem~211_combout ),
	.cout());
defparam \mem~211 .lut_mask = 16'hFFFE;
defparam \mem~211 .sum_lutc_input = "datac";

dffeas \mem~112 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~112_q ),
	.prn(vcc));
defparam \mem~112 .is_wysiwyg = "true";
defparam \mem~112 .power_up = "low";

cycloneive_lcell_comb \mem~129 (
	.dataa(\mem~80_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~128_combout ),
	.datad(\mem~112_q ),
	.cin(gnd),
	.combout(\mem~129_combout ),
	.cout());
defparam \mem~129 .lut_mask = 16'hFFBE;
defparam \mem~129 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~212 (
	.dataa(\wr_ptr[1]~q ),
	.datab(\write~combout ),
	.datac(\wr_ptr[2]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem~212_combout ),
	.cout());
defparam \mem~212 .lut_mask = 16'hEFFF;
defparam \mem~212 .sum_lutc_input = "datac";

dffeas \mem~32 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~32_q ),
	.prn(vcc));
defparam \mem~32 .is_wysiwyg = "true";
defparam \mem~32 .power_up = "low";

cycloneive_lcell_comb \mem~213 (
	.dataa(\wr_ptr[0]~q ),
	.datab(\write~combout ),
	.datac(\wr_ptr[2]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~213_combout ),
	.cout());
defparam \mem~213 .lut_mask = 16'hEFFF;
defparam \mem~213 .sum_lutc_input = "datac";

dffeas \mem~16 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~16_q ),
	.prn(vcc));
defparam \mem~16 .is_wysiwyg = "true";
defparam \mem~16 .power_up = "low";

cycloneive_lcell_comb \mem~214 (
	.dataa(\write~combout ),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~214_combout ),
	.cout());
defparam \mem~214 .lut_mask = 16'hBFFF;
defparam \mem~214 .sum_lutc_input = "datac";

dffeas \mem~0 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~0_q ),
	.prn(vcc));
defparam \mem~0 .is_wysiwyg = "true";
defparam \mem~0 .power_up = "low";

cycloneive_lcell_comb \mem~130 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~16_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~0_q ),
	.cin(gnd),
	.combout(\mem~130_combout ),
	.cout());
defparam \mem~130 .lut_mask = 16'hFFDE;
defparam \mem~130 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~215 (
	.dataa(\wr_ptr[0]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\write~combout ),
	.datad(\wr_ptr[2]~q ),
	.cin(gnd),
	.combout(\mem~215_combout ),
	.cout());
defparam \mem~215 .lut_mask = 16'hFEFF;
defparam \mem~215 .sum_lutc_input = "datac";

dffeas \mem~48 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~48_q ),
	.prn(vcc));
defparam \mem~48 .is_wysiwyg = "true";
defparam \mem~48 .power_up = "low";

cycloneive_lcell_comb \mem~131 (
	.dataa(\mem~32_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~130_combout ),
	.datad(\mem~48_q ),
	.cin(gnd),
	.combout(\mem~131_combout ),
	.cout());
defparam \mem~131 .lut_mask = 16'hFFBE;
defparam \mem~131 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~132 (
	.dataa(\mem~129_combout ),
	.datab(\mem~131_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~132_combout ),
	.cout());
defparam \mem~132 .lut_mask = 16'hAACC;
defparam \mem~132 .sum_lutc_input = "datac";

dffeas \internal_out_payload[0] (
	.clk(clk),
	.d(\mem~132_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[0]~q ),
	.prn(vcc));
defparam \internal_out_payload[0] .is_wysiwyg = "true";
defparam \internal_out_payload[0] .power_up = "low";

dffeas \mem~81 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~81_q ),
	.prn(vcc));
defparam \mem~81 .is_wysiwyg = "true";
defparam \mem~81 .power_up = "low";

dffeas \mem~97 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~97_q ),
	.prn(vcc));
defparam \mem~97 .is_wysiwyg = "true";
defparam \mem~97 .power_up = "low";

dffeas \mem~65 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~65_q ),
	.prn(vcc));
defparam \mem~65 .is_wysiwyg = "true";
defparam \mem~65 .power_up = "low";

cycloneive_lcell_comb \mem~133 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~97_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~65_q ),
	.cin(gnd),
	.combout(\mem~133_combout ),
	.cout());
defparam \mem~133 .lut_mask = 16'hFFDE;
defparam \mem~133 .sum_lutc_input = "datac";

dffeas \mem~113 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~113_q ),
	.prn(vcc));
defparam \mem~113 .is_wysiwyg = "true";
defparam \mem~113 .power_up = "low";

cycloneive_lcell_comb \mem~134 (
	.dataa(\mem~81_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~133_combout ),
	.datad(\mem~113_q ),
	.cin(gnd),
	.combout(\mem~134_combout ),
	.cout());
defparam \mem~134 .lut_mask = 16'hFFBE;
defparam \mem~134 .sum_lutc_input = "datac";

dffeas \mem~33 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~33_q ),
	.prn(vcc));
defparam \mem~33 .is_wysiwyg = "true";
defparam \mem~33 .power_up = "low";

dffeas \mem~17 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~17_q ),
	.prn(vcc));
defparam \mem~17 .is_wysiwyg = "true";
defparam \mem~17 .power_up = "low";

dffeas \mem~1 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~1_q ),
	.prn(vcc));
defparam \mem~1 .is_wysiwyg = "true";
defparam \mem~1 .power_up = "low";

cycloneive_lcell_comb \mem~135 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~17_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~1_q ),
	.cin(gnd),
	.combout(\mem~135_combout ),
	.cout());
defparam \mem~135 .lut_mask = 16'hFFDE;
defparam \mem~135 .sum_lutc_input = "datac";

dffeas \mem~49 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~49_q ),
	.prn(vcc));
defparam \mem~49 .is_wysiwyg = "true";
defparam \mem~49 .power_up = "low";

cycloneive_lcell_comb \mem~136 (
	.dataa(\mem~33_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~135_combout ),
	.datad(\mem~49_q ),
	.cin(gnd),
	.combout(\mem~136_combout ),
	.cout());
defparam \mem~136 .lut_mask = 16'hFFBE;
defparam \mem~136 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~137 (
	.dataa(\mem~134_combout ),
	.datab(\mem~136_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~137_combout ),
	.cout());
defparam \mem~137 .lut_mask = 16'hAACC;
defparam \mem~137 .sum_lutc_input = "datac";

dffeas \internal_out_payload[1] (
	.clk(clk),
	.d(\mem~137_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[1]~q ),
	.prn(vcc));
defparam \internal_out_payload[1] .is_wysiwyg = "true";
defparam \internal_out_payload[1] .power_up = "low";

dffeas \mem~82 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~82_q ),
	.prn(vcc));
defparam \mem~82 .is_wysiwyg = "true";
defparam \mem~82 .power_up = "low";

dffeas \mem~98 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~98_q ),
	.prn(vcc));
defparam \mem~98 .is_wysiwyg = "true";
defparam \mem~98 .power_up = "low";

dffeas \mem~66 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~66_q ),
	.prn(vcc));
defparam \mem~66 .is_wysiwyg = "true";
defparam \mem~66 .power_up = "low";

cycloneive_lcell_comb \mem~138 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~98_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~66_q ),
	.cin(gnd),
	.combout(\mem~138_combout ),
	.cout());
defparam \mem~138 .lut_mask = 16'hFFDE;
defparam \mem~138 .sum_lutc_input = "datac";

dffeas \mem~114 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~114_q ),
	.prn(vcc));
defparam \mem~114 .is_wysiwyg = "true";
defparam \mem~114 .power_up = "low";

cycloneive_lcell_comb \mem~139 (
	.dataa(\mem~82_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~138_combout ),
	.datad(\mem~114_q ),
	.cin(gnd),
	.combout(\mem~139_combout ),
	.cout());
defparam \mem~139 .lut_mask = 16'hFFBE;
defparam \mem~139 .sum_lutc_input = "datac";

dffeas \mem~34 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~34_q ),
	.prn(vcc));
defparam \mem~34 .is_wysiwyg = "true";
defparam \mem~34 .power_up = "low";

dffeas \mem~18 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~18_q ),
	.prn(vcc));
defparam \mem~18 .is_wysiwyg = "true";
defparam \mem~18 .power_up = "low";

dffeas \mem~2 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~2_q ),
	.prn(vcc));
defparam \mem~2 .is_wysiwyg = "true";
defparam \mem~2 .power_up = "low";

cycloneive_lcell_comb \mem~140 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~18_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~2_q ),
	.cin(gnd),
	.combout(\mem~140_combout ),
	.cout());
defparam \mem~140 .lut_mask = 16'hFFDE;
defparam \mem~140 .sum_lutc_input = "datac";

dffeas \mem~50 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~50_q ),
	.prn(vcc));
defparam \mem~50 .is_wysiwyg = "true";
defparam \mem~50 .power_up = "low";

cycloneive_lcell_comb \mem~141 (
	.dataa(\mem~34_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~140_combout ),
	.datad(\mem~50_q ),
	.cin(gnd),
	.combout(\mem~141_combout ),
	.cout());
defparam \mem~141 .lut_mask = 16'hFFBE;
defparam \mem~141 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~142 (
	.dataa(\mem~139_combout ),
	.datab(\mem~141_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~142_combout ),
	.cout());
defparam \mem~142 .lut_mask = 16'hAACC;
defparam \mem~142 .sum_lutc_input = "datac";

dffeas \internal_out_payload[2] (
	.clk(clk),
	.d(\mem~142_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[2]~q ),
	.prn(vcc));
defparam \internal_out_payload[2] .is_wysiwyg = "true";
defparam \internal_out_payload[2] .power_up = "low";

dffeas \mem~83 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~83_q ),
	.prn(vcc));
defparam \mem~83 .is_wysiwyg = "true";
defparam \mem~83 .power_up = "low";

dffeas \mem~99 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~99_q ),
	.prn(vcc));
defparam \mem~99 .is_wysiwyg = "true";
defparam \mem~99 .power_up = "low";

dffeas \mem~67 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~67_q ),
	.prn(vcc));
defparam \mem~67 .is_wysiwyg = "true";
defparam \mem~67 .power_up = "low";

cycloneive_lcell_comb \mem~143 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~99_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~67_q ),
	.cin(gnd),
	.combout(\mem~143_combout ),
	.cout());
defparam \mem~143 .lut_mask = 16'hFFDE;
defparam \mem~143 .sum_lutc_input = "datac";

dffeas \mem~115 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~115_q ),
	.prn(vcc));
defparam \mem~115 .is_wysiwyg = "true";
defparam \mem~115 .power_up = "low";

cycloneive_lcell_comb \mem~144 (
	.dataa(\mem~83_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~143_combout ),
	.datad(\mem~115_q ),
	.cin(gnd),
	.combout(\mem~144_combout ),
	.cout());
defparam \mem~144 .lut_mask = 16'hFFBE;
defparam \mem~144 .sum_lutc_input = "datac";

dffeas \mem~35 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~35_q ),
	.prn(vcc));
defparam \mem~35 .is_wysiwyg = "true";
defparam \mem~35 .power_up = "low";

dffeas \mem~19 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~19_q ),
	.prn(vcc));
defparam \mem~19 .is_wysiwyg = "true";
defparam \mem~19 .power_up = "low";

dffeas \mem~3 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~3_q ),
	.prn(vcc));
defparam \mem~3 .is_wysiwyg = "true";
defparam \mem~3 .power_up = "low";

cycloneive_lcell_comb \mem~145 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~19_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~3_q ),
	.cin(gnd),
	.combout(\mem~145_combout ),
	.cout());
defparam \mem~145 .lut_mask = 16'hFFDE;
defparam \mem~145 .sum_lutc_input = "datac";

dffeas \mem~51 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~51_q ),
	.prn(vcc));
defparam \mem~51 .is_wysiwyg = "true";
defparam \mem~51 .power_up = "low";

cycloneive_lcell_comb \mem~146 (
	.dataa(\mem~35_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~145_combout ),
	.datad(\mem~51_q ),
	.cin(gnd),
	.combout(\mem~146_combout ),
	.cout());
defparam \mem~146 .lut_mask = 16'hFFBE;
defparam \mem~146 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~147 (
	.dataa(\mem~144_combout ),
	.datab(\mem~146_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~147_combout ),
	.cout());
defparam \mem~147 .lut_mask = 16'hAACC;
defparam \mem~147 .sum_lutc_input = "datac";

dffeas \internal_out_payload[3] (
	.clk(clk),
	.d(\mem~147_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[3]~q ),
	.prn(vcc));
defparam \internal_out_payload[3] .is_wysiwyg = "true";
defparam \internal_out_payload[3] .power_up = "low";

dffeas \mem~84 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~84_q ),
	.prn(vcc));
defparam \mem~84 .is_wysiwyg = "true";
defparam \mem~84 .power_up = "low";

dffeas \mem~100 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~100_q ),
	.prn(vcc));
defparam \mem~100 .is_wysiwyg = "true";
defparam \mem~100 .power_up = "low";

dffeas \mem~68 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~68_q ),
	.prn(vcc));
defparam \mem~68 .is_wysiwyg = "true";
defparam \mem~68 .power_up = "low";

cycloneive_lcell_comb \mem~148 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~100_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~68_q ),
	.cin(gnd),
	.combout(\mem~148_combout ),
	.cout());
defparam \mem~148 .lut_mask = 16'hFFDE;
defparam \mem~148 .sum_lutc_input = "datac";

dffeas \mem~116 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~116_q ),
	.prn(vcc));
defparam \mem~116 .is_wysiwyg = "true";
defparam \mem~116 .power_up = "low";

cycloneive_lcell_comb \mem~149 (
	.dataa(\mem~84_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~148_combout ),
	.datad(\mem~116_q ),
	.cin(gnd),
	.combout(\mem~149_combout ),
	.cout());
defparam \mem~149 .lut_mask = 16'hFFBE;
defparam \mem~149 .sum_lutc_input = "datac";

dffeas \mem~36 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~36_q ),
	.prn(vcc));
defparam \mem~36 .is_wysiwyg = "true";
defparam \mem~36 .power_up = "low";

dffeas \mem~20 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~20_q ),
	.prn(vcc));
defparam \mem~20 .is_wysiwyg = "true";
defparam \mem~20 .power_up = "low";

dffeas \mem~4 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~4_q ),
	.prn(vcc));
defparam \mem~4 .is_wysiwyg = "true";
defparam \mem~4 .power_up = "low";

cycloneive_lcell_comb \mem~150 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~20_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~4_q ),
	.cin(gnd),
	.combout(\mem~150_combout ),
	.cout());
defparam \mem~150 .lut_mask = 16'hFFDE;
defparam \mem~150 .sum_lutc_input = "datac";

dffeas \mem~52 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~52_q ),
	.prn(vcc));
defparam \mem~52 .is_wysiwyg = "true";
defparam \mem~52 .power_up = "low";

cycloneive_lcell_comb \mem~151 (
	.dataa(\mem~36_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~150_combout ),
	.datad(\mem~52_q ),
	.cin(gnd),
	.combout(\mem~151_combout ),
	.cout());
defparam \mem~151 .lut_mask = 16'hFFBE;
defparam \mem~151 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~152 (
	.dataa(\mem~149_combout ),
	.datab(\mem~151_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~152_combout ),
	.cout());
defparam \mem~152 .lut_mask = 16'hAACC;
defparam \mem~152 .sum_lutc_input = "datac";

dffeas \internal_out_payload[4] (
	.clk(clk),
	.d(\mem~152_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[4]~q ),
	.prn(vcc));
defparam \internal_out_payload[4] .is_wysiwyg = "true";
defparam \internal_out_payload[4] .power_up = "low";

dffeas \mem~91 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~91_q ),
	.prn(vcc));
defparam \mem~91 .is_wysiwyg = "true";
defparam \mem~91 .power_up = "low";

dffeas \mem~107 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~107_q ),
	.prn(vcc));
defparam \mem~107 .is_wysiwyg = "true";
defparam \mem~107 .power_up = "low";

dffeas \mem~75 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~75_q ),
	.prn(vcc));
defparam \mem~75 .is_wysiwyg = "true";
defparam \mem~75 .power_up = "low";

cycloneive_lcell_comb \mem~153 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~107_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~75_q ),
	.cin(gnd),
	.combout(\mem~153_combout ),
	.cout());
defparam \mem~153 .lut_mask = 16'hFFDE;
defparam \mem~153 .sum_lutc_input = "datac";

dffeas \mem~123 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~123_q ),
	.prn(vcc));
defparam \mem~123 .is_wysiwyg = "true";
defparam \mem~123 .power_up = "low";

cycloneive_lcell_comb \mem~154 (
	.dataa(\mem~91_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~153_combout ),
	.datad(\mem~123_q ),
	.cin(gnd),
	.combout(\mem~154_combout ),
	.cout());
defparam \mem~154 .lut_mask = 16'hFFBE;
defparam \mem~154 .sum_lutc_input = "datac";

dffeas \mem~43 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~43_q ),
	.prn(vcc));
defparam \mem~43 .is_wysiwyg = "true";
defparam \mem~43 .power_up = "low";

dffeas \mem~27 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~27_q ),
	.prn(vcc));
defparam \mem~27 .is_wysiwyg = "true";
defparam \mem~27 .power_up = "low";

dffeas \mem~11 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~11_q ),
	.prn(vcc));
defparam \mem~11 .is_wysiwyg = "true";
defparam \mem~11 .power_up = "low";

cycloneive_lcell_comb \mem~155 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~27_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~11_q ),
	.cin(gnd),
	.combout(\mem~155_combout ),
	.cout());
defparam \mem~155 .lut_mask = 16'hFFDE;
defparam \mem~155 .sum_lutc_input = "datac";

dffeas \mem~59 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~59_q ),
	.prn(vcc));
defparam \mem~59 .is_wysiwyg = "true";
defparam \mem~59 .power_up = "low";

cycloneive_lcell_comb \mem~156 (
	.dataa(\mem~43_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~155_combout ),
	.datad(\mem~59_q ),
	.cin(gnd),
	.combout(\mem~156_combout ),
	.cout());
defparam \mem~156 .lut_mask = 16'hFFBE;
defparam \mem~156 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~157 (
	.dataa(\mem~154_combout ),
	.datab(\mem~156_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~157_combout ),
	.cout());
defparam \mem~157 .lut_mask = 16'hAACC;
defparam \mem~157 .sum_lutc_input = "datac";

dffeas \internal_out_payload[11] (
	.clk(clk),
	.d(\mem~157_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[11]~q ),
	.prn(vcc));
defparam \internal_out_payload[11] .is_wysiwyg = "true";
defparam \internal_out_payload[11] .power_up = "low";

dffeas \mem~93 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~93_q ),
	.prn(vcc));
defparam \mem~93 .is_wysiwyg = "true";
defparam \mem~93 .power_up = "low";

dffeas \mem~109 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~109_q ),
	.prn(vcc));
defparam \mem~109 .is_wysiwyg = "true";
defparam \mem~109 .power_up = "low";

dffeas \mem~77 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~77_q ),
	.prn(vcc));
defparam \mem~77 .is_wysiwyg = "true";
defparam \mem~77 .power_up = "low";

cycloneive_lcell_comb \mem~158 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~109_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~77_q ),
	.cin(gnd),
	.combout(\mem~158_combout ),
	.cout());
defparam \mem~158 .lut_mask = 16'hFFDE;
defparam \mem~158 .sum_lutc_input = "datac";

dffeas \mem~125 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~125_q ),
	.prn(vcc));
defparam \mem~125 .is_wysiwyg = "true";
defparam \mem~125 .power_up = "low";

cycloneive_lcell_comb \mem~159 (
	.dataa(\mem~93_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~158_combout ),
	.datad(\mem~125_q ),
	.cin(gnd),
	.combout(\mem~159_combout ),
	.cout());
defparam \mem~159 .lut_mask = 16'hFFBE;
defparam \mem~159 .sum_lutc_input = "datac";

dffeas \mem~45 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~45_q ),
	.prn(vcc));
defparam \mem~45 .is_wysiwyg = "true";
defparam \mem~45 .power_up = "low";

dffeas \mem~29 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~29_q ),
	.prn(vcc));
defparam \mem~29 .is_wysiwyg = "true";
defparam \mem~29 .power_up = "low";

dffeas \mem~13 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~13_q ),
	.prn(vcc));
defparam \mem~13 .is_wysiwyg = "true";
defparam \mem~13 .power_up = "low";

cycloneive_lcell_comb \mem~160 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~29_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~13_q ),
	.cin(gnd),
	.combout(\mem~160_combout ),
	.cout());
defparam \mem~160 .lut_mask = 16'hFFDE;
defparam \mem~160 .sum_lutc_input = "datac";

dffeas \mem~61 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~61_q ),
	.prn(vcc));
defparam \mem~61 .is_wysiwyg = "true";
defparam \mem~61 .power_up = "low";

cycloneive_lcell_comb \mem~161 (
	.dataa(\mem~45_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~160_combout ),
	.datad(\mem~61_q ),
	.cin(gnd),
	.combout(\mem~161_combout ),
	.cout());
defparam \mem~161 .lut_mask = 16'hFFBE;
defparam \mem~161 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~162 (
	.dataa(\mem~159_combout ),
	.datab(\mem~161_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~162_combout ),
	.cout());
defparam \mem~162 .lut_mask = 16'hAACC;
defparam \mem~162 .sum_lutc_input = "datac";

dffeas \internal_out_payload[13] (
	.clk(clk),
	.d(\mem~162_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[13]~q ),
	.prn(vcc));
defparam \internal_out_payload[13] .is_wysiwyg = "true";
defparam \internal_out_payload[13] .power_up = "low";

dffeas \mem~92 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~92_q ),
	.prn(vcc));
defparam \mem~92 .is_wysiwyg = "true";
defparam \mem~92 .power_up = "low";

dffeas \mem~108 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~108_q ),
	.prn(vcc));
defparam \mem~108 .is_wysiwyg = "true";
defparam \mem~108 .power_up = "low";

dffeas \mem~76 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~76_q ),
	.prn(vcc));
defparam \mem~76 .is_wysiwyg = "true";
defparam \mem~76 .power_up = "low";

cycloneive_lcell_comb \mem~163 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~108_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~76_q ),
	.cin(gnd),
	.combout(\mem~163_combout ),
	.cout());
defparam \mem~163 .lut_mask = 16'hFFDE;
defparam \mem~163 .sum_lutc_input = "datac";

dffeas \mem~124 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~124_q ),
	.prn(vcc));
defparam \mem~124 .is_wysiwyg = "true";
defparam \mem~124 .power_up = "low";

cycloneive_lcell_comb \mem~164 (
	.dataa(\mem~92_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~163_combout ),
	.datad(\mem~124_q ),
	.cin(gnd),
	.combout(\mem~164_combout ),
	.cout());
defparam \mem~164 .lut_mask = 16'hFFBE;
defparam \mem~164 .sum_lutc_input = "datac";

dffeas \mem~44 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~44_q ),
	.prn(vcc));
defparam \mem~44 .is_wysiwyg = "true";
defparam \mem~44 .power_up = "low";

dffeas \mem~28 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~28_q ),
	.prn(vcc));
defparam \mem~28 .is_wysiwyg = "true";
defparam \mem~28 .power_up = "low";

dffeas \mem~12 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~12_q ),
	.prn(vcc));
defparam \mem~12 .is_wysiwyg = "true";
defparam \mem~12 .power_up = "low";

cycloneive_lcell_comb \mem~165 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~28_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~12_q ),
	.cin(gnd),
	.combout(\mem~165_combout ),
	.cout());
defparam \mem~165 .lut_mask = 16'hFFDE;
defparam \mem~165 .sum_lutc_input = "datac";

dffeas \mem~60 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~60_q ),
	.prn(vcc));
defparam \mem~60 .is_wysiwyg = "true";
defparam \mem~60 .power_up = "low";

cycloneive_lcell_comb \mem~166 (
	.dataa(\mem~44_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~165_combout ),
	.datad(\mem~60_q ),
	.cin(gnd),
	.combout(\mem~166_combout ),
	.cout());
defparam \mem~166 .lut_mask = 16'hFFBE;
defparam \mem~166 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~167 (
	.dataa(\mem~164_combout ),
	.datab(\mem~166_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~167_combout ),
	.cout());
defparam \mem~167 .lut_mask = 16'hAACC;
defparam \mem~167 .sum_lutc_input = "datac";

dffeas \internal_out_payload[12] (
	.clk(clk),
	.d(\mem~167_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[12]~q ),
	.prn(vcc));
defparam \internal_out_payload[12] .is_wysiwyg = "true";
defparam \internal_out_payload[12] .power_up = "low";

dffeas \mem~85 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~85_q ),
	.prn(vcc));
defparam \mem~85 .is_wysiwyg = "true";
defparam \mem~85 .power_up = "low";

dffeas \mem~101 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~101_q ),
	.prn(vcc));
defparam \mem~101 .is_wysiwyg = "true";
defparam \mem~101 .power_up = "low";

dffeas \mem~69 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~69_q ),
	.prn(vcc));
defparam \mem~69 .is_wysiwyg = "true";
defparam \mem~69 .power_up = "low";

cycloneive_lcell_comb \mem~168 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~101_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~69_q ),
	.cin(gnd),
	.combout(\mem~168_combout ),
	.cout());
defparam \mem~168 .lut_mask = 16'hFFDE;
defparam \mem~168 .sum_lutc_input = "datac";

dffeas \mem~117 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~117_q ),
	.prn(vcc));
defparam \mem~117 .is_wysiwyg = "true";
defparam \mem~117 .power_up = "low";

cycloneive_lcell_comb \mem~169 (
	.dataa(\mem~85_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~168_combout ),
	.datad(\mem~117_q ),
	.cin(gnd),
	.combout(\mem~169_combout ),
	.cout());
defparam \mem~169 .lut_mask = 16'hFFBE;
defparam \mem~169 .sum_lutc_input = "datac";

dffeas \mem~37 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~37_q ),
	.prn(vcc));
defparam \mem~37 .is_wysiwyg = "true";
defparam \mem~37 .power_up = "low";

dffeas \mem~21 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~21_q ),
	.prn(vcc));
defparam \mem~21 .is_wysiwyg = "true";
defparam \mem~21 .power_up = "low";

dffeas \mem~5 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~5_q ),
	.prn(vcc));
defparam \mem~5 .is_wysiwyg = "true";
defparam \mem~5 .power_up = "low";

cycloneive_lcell_comb \mem~170 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~21_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~5_q ),
	.cin(gnd),
	.combout(\mem~170_combout ),
	.cout());
defparam \mem~170 .lut_mask = 16'hFFDE;
defparam \mem~170 .sum_lutc_input = "datac";

dffeas \mem~53 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~53_q ),
	.prn(vcc));
defparam \mem~53 .is_wysiwyg = "true";
defparam \mem~53 .power_up = "low";

cycloneive_lcell_comb \mem~171 (
	.dataa(\mem~37_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~170_combout ),
	.datad(\mem~53_q ),
	.cin(gnd),
	.combout(\mem~171_combout ),
	.cout());
defparam \mem~171 .lut_mask = 16'hFFBE;
defparam \mem~171 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~172 (
	.dataa(\mem~169_combout ),
	.datab(\mem~171_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~172_combout ),
	.cout());
defparam \mem~172 .lut_mask = 16'hAACC;
defparam \mem~172 .sum_lutc_input = "datac";

dffeas \internal_out_payload[5] (
	.clk(clk),
	.d(\mem~172_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[5]~q ),
	.prn(vcc));
defparam \internal_out_payload[5] .is_wysiwyg = "true";
defparam \internal_out_payload[5] .power_up = "low";

dffeas \mem~94 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~94_q ),
	.prn(vcc));
defparam \mem~94 .is_wysiwyg = "true";
defparam \mem~94 .power_up = "low";

dffeas \mem~110 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~110_q ),
	.prn(vcc));
defparam \mem~110 .is_wysiwyg = "true";
defparam \mem~110 .power_up = "low";

dffeas \mem~78 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~78_q ),
	.prn(vcc));
defparam \mem~78 .is_wysiwyg = "true";
defparam \mem~78 .power_up = "low";

cycloneive_lcell_comb \mem~173 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~110_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~78_q ),
	.cin(gnd),
	.combout(\mem~173_combout ),
	.cout());
defparam \mem~173 .lut_mask = 16'hFFDE;
defparam \mem~173 .sum_lutc_input = "datac";

dffeas \mem~126 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~126_q ),
	.prn(vcc));
defparam \mem~126 .is_wysiwyg = "true";
defparam \mem~126 .power_up = "low";

cycloneive_lcell_comb \mem~174 (
	.dataa(\mem~94_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~173_combout ),
	.datad(\mem~126_q ),
	.cin(gnd),
	.combout(\mem~174_combout ),
	.cout());
defparam \mem~174 .lut_mask = 16'hFFBE;
defparam \mem~174 .sum_lutc_input = "datac";

dffeas \mem~46 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~46_q ),
	.prn(vcc));
defparam \mem~46 .is_wysiwyg = "true";
defparam \mem~46 .power_up = "low";

dffeas \mem~30 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~30_q ),
	.prn(vcc));
defparam \mem~30 .is_wysiwyg = "true";
defparam \mem~30 .power_up = "low";

dffeas \mem~14 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~14_q ),
	.prn(vcc));
defparam \mem~14 .is_wysiwyg = "true";
defparam \mem~14 .power_up = "low";

cycloneive_lcell_comb \mem~175 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~30_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~14_q ),
	.cin(gnd),
	.combout(\mem~175_combout ),
	.cout());
defparam \mem~175 .lut_mask = 16'hFFDE;
defparam \mem~175 .sum_lutc_input = "datac";

dffeas \mem~62 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~62_q ),
	.prn(vcc));
defparam \mem~62 .is_wysiwyg = "true";
defparam \mem~62 .power_up = "low";

cycloneive_lcell_comb \mem~176 (
	.dataa(\mem~46_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~175_combout ),
	.datad(\mem~62_q ),
	.cin(gnd),
	.combout(\mem~176_combout ),
	.cout());
defparam \mem~176 .lut_mask = 16'hFFBE;
defparam \mem~176 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~177 (
	.dataa(\mem~174_combout ),
	.datab(\mem~176_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~177_combout ),
	.cout());
defparam \mem~177 .lut_mask = 16'hAACC;
defparam \mem~177 .sum_lutc_input = "datac";

dffeas \internal_out_payload[14] (
	.clk(clk),
	.d(\mem~177_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[14]~q ),
	.prn(vcc));
defparam \internal_out_payload[14] .is_wysiwyg = "true";
defparam \internal_out_payload[14] .power_up = "low";

dffeas \mem~95 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~95_q ),
	.prn(vcc));
defparam \mem~95 .is_wysiwyg = "true";
defparam \mem~95 .power_up = "low";

dffeas \mem~111 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~111_q ),
	.prn(vcc));
defparam \mem~111 .is_wysiwyg = "true";
defparam \mem~111 .power_up = "low";

dffeas \mem~79 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~79_q ),
	.prn(vcc));
defparam \mem~79 .is_wysiwyg = "true";
defparam \mem~79 .power_up = "low";

cycloneive_lcell_comb \mem~178 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~111_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~79_q ),
	.cin(gnd),
	.combout(\mem~178_combout ),
	.cout());
defparam \mem~178 .lut_mask = 16'hFFDE;
defparam \mem~178 .sum_lutc_input = "datac";

dffeas \mem~127 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~127_q ),
	.prn(vcc));
defparam \mem~127 .is_wysiwyg = "true";
defparam \mem~127 .power_up = "low";

cycloneive_lcell_comb \mem~179 (
	.dataa(\mem~95_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~178_combout ),
	.datad(\mem~127_q ),
	.cin(gnd),
	.combout(\mem~179_combout ),
	.cout());
defparam \mem~179 .lut_mask = 16'hFFBE;
defparam \mem~179 .sum_lutc_input = "datac";

dffeas \mem~47 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~47_q ),
	.prn(vcc));
defparam \mem~47 .is_wysiwyg = "true";
defparam \mem~47 .power_up = "low";

dffeas \mem~31 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~31_q ),
	.prn(vcc));
defparam \mem~31 .is_wysiwyg = "true";
defparam \mem~31 .power_up = "low";

dffeas \mem~15 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~15_q ),
	.prn(vcc));
defparam \mem~15 .is_wysiwyg = "true";
defparam \mem~15 .power_up = "low";

cycloneive_lcell_comb \mem~180 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~31_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~15_q ),
	.cin(gnd),
	.combout(\mem~180_combout ),
	.cout());
defparam \mem~180 .lut_mask = 16'hFFDE;
defparam \mem~180 .sum_lutc_input = "datac";

dffeas \mem~63 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~63_q ),
	.prn(vcc));
defparam \mem~63 .is_wysiwyg = "true";
defparam \mem~63 .power_up = "low";

cycloneive_lcell_comb \mem~181 (
	.dataa(\mem~47_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~180_combout ),
	.datad(\mem~63_q ),
	.cin(gnd),
	.combout(\mem~181_combout ),
	.cout());
defparam \mem~181 .lut_mask = 16'hFFBE;
defparam \mem~181 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~182 (
	.dataa(\mem~179_combout ),
	.datab(\mem~181_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~182_combout ),
	.cout());
defparam \mem~182 .lut_mask = 16'hAACC;
defparam \mem~182 .sum_lutc_input = "datac";

dffeas \internal_out_payload[15] (
	.clk(clk),
	.d(\mem~182_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[15]~q ),
	.prn(vcc));
defparam \internal_out_payload[15] .is_wysiwyg = "true";
defparam \internal_out_payload[15] .power_up = "low";

dffeas \mem~90 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~90_q ),
	.prn(vcc));
defparam \mem~90 .is_wysiwyg = "true";
defparam \mem~90 .power_up = "low";

dffeas \mem~106 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~106_q ),
	.prn(vcc));
defparam \mem~106 .is_wysiwyg = "true";
defparam \mem~106 .power_up = "low";

dffeas \mem~74 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~74_q ),
	.prn(vcc));
defparam \mem~74 .is_wysiwyg = "true";
defparam \mem~74 .power_up = "low";

cycloneive_lcell_comb \mem~183 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~106_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~74_q ),
	.cin(gnd),
	.combout(\mem~183_combout ),
	.cout());
defparam \mem~183 .lut_mask = 16'hFFDE;
defparam \mem~183 .sum_lutc_input = "datac";

dffeas \mem~122 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~122_q ),
	.prn(vcc));
defparam \mem~122 .is_wysiwyg = "true";
defparam \mem~122 .power_up = "low";

cycloneive_lcell_comb \mem~184 (
	.dataa(\mem~90_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~183_combout ),
	.datad(\mem~122_q ),
	.cin(gnd),
	.combout(\mem~184_combout ),
	.cout());
defparam \mem~184 .lut_mask = 16'hFFBE;
defparam \mem~184 .sum_lutc_input = "datac";

dffeas \mem~42 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~42_q ),
	.prn(vcc));
defparam \mem~42 .is_wysiwyg = "true";
defparam \mem~42 .power_up = "low";

dffeas \mem~26 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~26_q ),
	.prn(vcc));
defparam \mem~26 .is_wysiwyg = "true";
defparam \mem~26 .power_up = "low";

dffeas \mem~10 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~10_q ),
	.prn(vcc));
defparam \mem~10 .is_wysiwyg = "true";
defparam \mem~10 .power_up = "low";

cycloneive_lcell_comb \mem~185 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~26_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~10_q ),
	.cin(gnd),
	.combout(\mem~185_combout ),
	.cout());
defparam \mem~185 .lut_mask = 16'hFFDE;
defparam \mem~185 .sum_lutc_input = "datac";

dffeas \mem~58 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~58_q ),
	.prn(vcc));
defparam \mem~58 .is_wysiwyg = "true";
defparam \mem~58 .power_up = "low";

cycloneive_lcell_comb \mem~186 (
	.dataa(\mem~42_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~185_combout ),
	.datad(\mem~58_q ),
	.cin(gnd),
	.combout(\mem~186_combout ),
	.cout());
defparam \mem~186 .lut_mask = 16'hFFBE;
defparam \mem~186 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~187 (
	.dataa(\mem~184_combout ),
	.datab(\mem~186_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~187_combout ),
	.cout());
defparam \mem~187 .lut_mask = 16'hAACC;
defparam \mem~187 .sum_lutc_input = "datac";

dffeas \internal_out_payload[10] (
	.clk(clk),
	.d(\mem~187_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[10]~q ),
	.prn(vcc));
defparam \internal_out_payload[10] .is_wysiwyg = "true";
defparam \internal_out_payload[10] .power_up = "low";

dffeas \mem~89 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~89_q ),
	.prn(vcc));
defparam \mem~89 .is_wysiwyg = "true";
defparam \mem~89 .power_up = "low";

dffeas \mem~105 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~105_q ),
	.prn(vcc));
defparam \mem~105 .is_wysiwyg = "true";
defparam \mem~105 .power_up = "low";

dffeas \mem~73 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~73_q ),
	.prn(vcc));
defparam \mem~73 .is_wysiwyg = "true";
defparam \mem~73 .power_up = "low";

cycloneive_lcell_comb \mem~188 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~105_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~73_q ),
	.cin(gnd),
	.combout(\mem~188_combout ),
	.cout());
defparam \mem~188 .lut_mask = 16'hFFDE;
defparam \mem~188 .sum_lutc_input = "datac";

dffeas \mem~121 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~121_q ),
	.prn(vcc));
defparam \mem~121 .is_wysiwyg = "true";
defparam \mem~121 .power_up = "low";

cycloneive_lcell_comb \mem~189 (
	.dataa(\mem~89_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~188_combout ),
	.datad(\mem~121_q ),
	.cin(gnd),
	.combout(\mem~189_combout ),
	.cout());
defparam \mem~189 .lut_mask = 16'hFFBE;
defparam \mem~189 .sum_lutc_input = "datac";

dffeas \mem~41 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~41_q ),
	.prn(vcc));
defparam \mem~41 .is_wysiwyg = "true";
defparam \mem~41 .power_up = "low";

dffeas \mem~25 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~25_q ),
	.prn(vcc));
defparam \mem~25 .is_wysiwyg = "true";
defparam \mem~25 .power_up = "low";

dffeas \mem~9 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~9_q ),
	.prn(vcc));
defparam \mem~9 .is_wysiwyg = "true";
defparam \mem~9 .power_up = "low";

cycloneive_lcell_comb \mem~190 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~25_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~9_q ),
	.cin(gnd),
	.combout(\mem~190_combout ),
	.cout());
defparam \mem~190 .lut_mask = 16'hFFDE;
defparam \mem~190 .sum_lutc_input = "datac";

dffeas \mem~57 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~57_q ),
	.prn(vcc));
defparam \mem~57 .is_wysiwyg = "true";
defparam \mem~57 .power_up = "low";

cycloneive_lcell_comb \mem~191 (
	.dataa(\mem~41_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~190_combout ),
	.datad(\mem~57_q ),
	.cin(gnd),
	.combout(\mem~191_combout ),
	.cout());
defparam \mem~191 .lut_mask = 16'hFFBE;
defparam \mem~191 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~192 (
	.dataa(\mem~189_combout ),
	.datab(\mem~191_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~192_combout ),
	.cout());
defparam \mem~192 .lut_mask = 16'hAACC;
defparam \mem~192 .sum_lutc_input = "datac";

dffeas \internal_out_payload[9] (
	.clk(clk),
	.d(\mem~192_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[9]~q ),
	.prn(vcc));
defparam \internal_out_payload[9] .is_wysiwyg = "true";
defparam \internal_out_payload[9] .power_up = "low";

dffeas \mem~88 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~88_q ),
	.prn(vcc));
defparam \mem~88 .is_wysiwyg = "true";
defparam \mem~88 .power_up = "low";

dffeas \mem~104 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~104_q ),
	.prn(vcc));
defparam \mem~104 .is_wysiwyg = "true";
defparam \mem~104 .power_up = "low";

dffeas \mem~72 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~72_q ),
	.prn(vcc));
defparam \mem~72 .is_wysiwyg = "true";
defparam \mem~72 .power_up = "low";

cycloneive_lcell_comb \mem~193 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~104_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~72_q ),
	.cin(gnd),
	.combout(\mem~193_combout ),
	.cout());
defparam \mem~193 .lut_mask = 16'hFFDE;
defparam \mem~193 .sum_lutc_input = "datac";

dffeas \mem~120 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~120_q ),
	.prn(vcc));
defparam \mem~120 .is_wysiwyg = "true";
defparam \mem~120 .power_up = "low";

cycloneive_lcell_comb \mem~194 (
	.dataa(\mem~88_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~193_combout ),
	.datad(\mem~120_q ),
	.cin(gnd),
	.combout(\mem~194_combout ),
	.cout());
defparam \mem~194 .lut_mask = 16'hFFBE;
defparam \mem~194 .sum_lutc_input = "datac";

dffeas \mem~40 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~40_q ),
	.prn(vcc));
defparam \mem~40 .is_wysiwyg = "true";
defparam \mem~40 .power_up = "low";

dffeas \mem~24 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~24_q ),
	.prn(vcc));
defparam \mem~24 .is_wysiwyg = "true";
defparam \mem~24 .power_up = "low";

dffeas \mem~8 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~8_q ),
	.prn(vcc));
defparam \mem~8 .is_wysiwyg = "true";
defparam \mem~8 .power_up = "low";

cycloneive_lcell_comb \mem~195 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~24_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~8_q ),
	.cin(gnd),
	.combout(\mem~195_combout ),
	.cout());
defparam \mem~195 .lut_mask = 16'hFFDE;
defparam \mem~195 .sum_lutc_input = "datac";

dffeas \mem~56 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~56_q ),
	.prn(vcc));
defparam \mem~56 .is_wysiwyg = "true";
defparam \mem~56 .power_up = "low";

cycloneive_lcell_comb \mem~196 (
	.dataa(\mem~40_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~195_combout ),
	.datad(\mem~56_q ),
	.cin(gnd),
	.combout(\mem~196_combout ),
	.cout());
defparam \mem~196 .lut_mask = 16'hFFBE;
defparam \mem~196 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~197 (
	.dataa(\mem~194_combout ),
	.datab(\mem~196_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~197_combout ),
	.cout());
defparam \mem~197 .lut_mask = 16'hAACC;
defparam \mem~197 .sum_lutc_input = "datac";

dffeas \internal_out_payload[8] (
	.clk(clk),
	.d(\mem~197_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[8]~q ),
	.prn(vcc));
defparam \internal_out_payload[8] .is_wysiwyg = "true";
defparam \internal_out_payload[8] .power_up = "low";

dffeas \mem~87 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~87_q ),
	.prn(vcc));
defparam \mem~87 .is_wysiwyg = "true";
defparam \mem~87 .power_up = "low";

dffeas \mem~103 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~103_q ),
	.prn(vcc));
defparam \mem~103 .is_wysiwyg = "true";
defparam \mem~103 .power_up = "low";

dffeas \mem~71 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~71_q ),
	.prn(vcc));
defparam \mem~71 .is_wysiwyg = "true";
defparam \mem~71 .power_up = "low";

cycloneive_lcell_comb \mem~198 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~103_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~71_q ),
	.cin(gnd),
	.combout(\mem~198_combout ),
	.cout());
defparam \mem~198 .lut_mask = 16'hFFDE;
defparam \mem~198 .sum_lutc_input = "datac";

dffeas \mem~119 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~119_q ),
	.prn(vcc));
defparam \mem~119 .is_wysiwyg = "true";
defparam \mem~119 .power_up = "low";

cycloneive_lcell_comb \mem~199 (
	.dataa(\mem~87_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~198_combout ),
	.datad(\mem~119_q ),
	.cin(gnd),
	.combout(\mem~199_combout ),
	.cout());
defparam \mem~199 .lut_mask = 16'hFFBE;
defparam \mem~199 .sum_lutc_input = "datac";

dffeas \mem~39 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~39_q ),
	.prn(vcc));
defparam \mem~39 .is_wysiwyg = "true";
defparam \mem~39 .power_up = "low";

dffeas \mem~23 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~23_q ),
	.prn(vcc));
defparam \mem~23 .is_wysiwyg = "true";
defparam \mem~23 .power_up = "low";

dffeas \mem~7 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~7_q ),
	.prn(vcc));
defparam \mem~7 .is_wysiwyg = "true";
defparam \mem~7 .power_up = "low";

cycloneive_lcell_comb \mem~200 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~23_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~7_q ),
	.cin(gnd),
	.combout(\mem~200_combout ),
	.cout());
defparam \mem~200 .lut_mask = 16'hFFDE;
defparam \mem~200 .sum_lutc_input = "datac";

dffeas \mem~55 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~55_q ),
	.prn(vcc));
defparam \mem~55 .is_wysiwyg = "true";
defparam \mem~55 .power_up = "low";

cycloneive_lcell_comb \mem~201 (
	.dataa(\mem~39_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~200_combout ),
	.datad(\mem~55_q ),
	.cin(gnd),
	.combout(\mem~201_combout ),
	.cout());
defparam \mem~201 .lut_mask = 16'hFFBE;
defparam \mem~201 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~202 (
	.dataa(\mem~199_combout ),
	.datab(\mem~201_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~202_combout ),
	.cout());
defparam \mem~202 .lut_mask = 16'hAACC;
defparam \mem~202 .sum_lutc_input = "datac";

dffeas \internal_out_payload[7] (
	.clk(clk),
	.d(\mem~202_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[7]~q ),
	.prn(vcc));
defparam \internal_out_payload[7] .is_wysiwyg = "true";
defparam \internal_out_payload[7] .power_up = "low";

dffeas \mem~86 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~208_combout ),
	.q(\mem~86_q ),
	.prn(vcc));
defparam \mem~86 .is_wysiwyg = "true";
defparam \mem~86 .power_up = "low";

dffeas \mem~102 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~209_combout ),
	.q(\mem~102_q ),
	.prn(vcc));
defparam \mem~102 .is_wysiwyg = "true";
defparam \mem~102 .power_up = "low";

dffeas \mem~70 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~210_combout ),
	.q(\mem~70_q ),
	.prn(vcc));
defparam \mem~70 .is_wysiwyg = "true";
defparam \mem~70 .power_up = "low";

cycloneive_lcell_comb \mem~203 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~102_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~70_q ),
	.cin(gnd),
	.combout(\mem~203_combout ),
	.cout());
defparam \mem~203 .lut_mask = 16'hFFDE;
defparam \mem~203 .sum_lutc_input = "datac";

dffeas \mem~118 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~211_combout ),
	.q(\mem~118_q ),
	.prn(vcc));
defparam \mem~118 .is_wysiwyg = "true";
defparam \mem~118 .power_up = "low";

cycloneive_lcell_comb \mem~204 (
	.dataa(\mem~86_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~203_combout ),
	.datad(\mem~118_q ),
	.cin(gnd),
	.combout(\mem~204_combout ),
	.cout());
defparam \mem~204 .lut_mask = 16'hFFBE;
defparam \mem~204 .sum_lutc_input = "datac";

dffeas \mem~38 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~212_combout ),
	.q(\mem~38_q ),
	.prn(vcc));
defparam \mem~38 .is_wysiwyg = "true";
defparam \mem~38 .power_up = "low";

dffeas \mem~22 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~213_combout ),
	.q(\mem~22_q ),
	.prn(vcc));
defparam \mem~22 .is_wysiwyg = "true";
defparam \mem~22 .power_up = "low";

dffeas \mem~6 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~214_combout ),
	.q(\mem~6_q ),
	.prn(vcc));
defparam \mem~6 .is_wysiwyg = "true";
defparam \mem~6 .power_up = "low";

cycloneive_lcell_comb \mem~205 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~22_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~6_q ),
	.cin(gnd),
	.combout(\mem~205_combout ),
	.cout());
defparam \mem~205 .lut_mask = 16'hFFDE;
defparam \mem~205 .sum_lutc_input = "datac";

dffeas \mem~54 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~215_combout ),
	.q(\mem~54_q ),
	.prn(vcc));
defparam \mem~54 .is_wysiwyg = "true";
defparam \mem~54 .power_up = "low";

cycloneive_lcell_comb \mem~206 (
	.dataa(\mem~38_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~205_combout ),
	.datad(\mem~54_q ),
	.cin(gnd),
	.combout(\mem~206_combout ),
	.cout());
defparam \mem~206 .lut_mask = 16'hFFBE;
defparam \mem~206 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~207 (
	.dataa(\mem~204_combout ),
	.datab(\mem~206_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~207_combout ),
	.cout());
defparam \mem~207 .lut_mask = 16'hAACC;
defparam \mem~207 .sum_lutc_input = "datac";

dffeas \internal_out_payload[6] (
	.clk(clk),
	.d(\mem~207_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[6]~q ),
	.prn(vcc));
defparam \internal_out_payload[6] .is_wysiwyg = "true";
defparam \internal_out_payload[6] .power_up = "low";

endmodule

module niosII_altera_avalon_sc_fifo_13 (
	clk,
	address_reg_1,
	reset,
	saved_grant_0,
	use_reg,
	saved_grant_1,
	WideOr1,
	mem_used_7,
	src_data_66,
	out_valid,
	mem_used_0,
	mem_87_0,
	mem_88_0,
	mem_54_0,
	mem_19_0,
	comb,
	mem_66_0,
	mem_48_0,
	out_endofpacket,
	mem_57_0,
	cp_ready,
	rf_source_data_87)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	address_reg_1;
input 	reset;
input 	saved_grant_0;
input 	use_reg;
input 	saved_grant_1;
input 	WideOr1;
output 	mem_used_7;
input 	src_data_66;
input 	out_valid;
output 	mem_used_0;
output 	mem_87_0;
output 	mem_88_0;
output 	mem_54_0;
output 	mem_19_0;
input 	comb;
output 	mem_66_0;
output 	mem_48_0;
input 	out_endofpacket;
output 	mem_57_0;
input 	cp_ready;
input 	rf_source_data_87;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used~6_combout ;
wire \mem_used[6]~4_combout ;
wire \mem_used[6]~5_combout ;
wire \mem_used[1]~q ;
wire \mem_used~8_combout ;
wire \mem_used[2]~q ;
wire \mem_used~10_combout ;
wire \mem_used[3]~q ;
wire \mem_used~9_combout ;
wire \mem_used[4]~q ;
wire \mem_used~7_combout ;
wire \mem_used[5]~q ;
wire \mem_used~3_combout ;
wire \mem_used[6]~q ;
wire \mem_used[7]~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem_used[0]~2_combout ;
wire \mem[7][87]~q ;
wire \mem~41_combout ;
wire \always6~0_combout ;
wire \mem[6][87]~q ;
wire \mem~34_combout ;
wire \always5~0_combout ;
wire \mem[5][87]~q ;
wire \mem~27_combout ;
wire \always4~0_combout ;
wire \mem[4][87]~q ;
wire \mem~20_combout ;
wire \always3~0_combout ;
wire \mem[3][87]~q ;
wire \mem~13_combout ;
wire \always2~0_combout ;
wire \mem[2][87]~q ;
wire \mem~6_combout ;
wire \always1~0_combout ;
wire \mem[1][87]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[7][88]~q ;
wire \mem~42_combout ;
wire \mem[6][88]~q ;
wire \mem~35_combout ;
wire \mem[5][88]~q ;
wire \mem~28_combout ;
wire \mem[4][88]~q ;
wire \mem~21_combout ;
wire \mem[3][88]~q ;
wire \mem~14_combout ;
wire \mem[2][88]~q ;
wire \mem~7_combout ;
wire \mem[1][88]~q ;
wire \mem~1_combout ;
wire \mem[7][85]~q ;
wire \mem~43_combout ;
wire \mem[6][54]~q ;
wire \mem~36_combout ;
wire \mem[5][54]~q ;
wire \mem~29_combout ;
wire \mem[4][54]~q ;
wire \mem~22_combout ;
wire \mem[3][54]~q ;
wire \mem~15_combout ;
wire \mem[2][54]~q ;
wire \mem~8_combout ;
wire \mem[1][54]~q ;
wire \mem~2_combout ;
wire \mem[7][19]~q ;
wire \mem~45_combout ;
wire \mem[6][19]~q ;
wire \mem~38_combout ;
wire \mem[5][19]~q ;
wire \mem~31_combout ;
wire \mem[4][19]~q ;
wire \mem~24_combout ;
wire \mem[3][19]~q ;
wire \mem~17_combout ;
wire \mem[2][19]~q ;
wire \mem~10_combout ;
wire \mem[1][19]~q ;
wire \mem~3_combout ;
wire \mem[7][66]~q ;
wire \mem~46_combout ;
wire \mem[6][66]~q ;
wire \mem~39_combout ;
wire \mem[5][66]~q ;
wire \mem~32_combout ;
wire \mem[4][66]~q ;
wire \mem~25_combout ;
wire \mem[3][66]~q ;
wire \mem~18_combout ;
wire \mem[2][66]~q ;
wire \mem~11_combout ;
wire \mem[1][66]~q ;
wire \mem~4_combout ;
wire \mem[7][48]~q ;
wire \mem~47_combout ;
wire \mem[6][48]~q ;
wire \mem~40_combout ;
wire \mem[5][48]~q ;
wire \mem~33_combout ;
wire \mem[4][48]~q ;
wire \mem~26_combout ;
wire \mem[3][48]~q ;
wire \mem~19_combout ;
wire \mem[2][48]~q ;
wire \mem~12_combout ;
wire \mem[1][48]~q ;
wire \mem~5_combout ;
wire \mem[7][57]~q ;
wire \mem~48_combout ;
wire \mem[6][57]~q ;
wire \mem~44_combout ;
wire \mem[5][57]~q ;
wire \mem~37_combout ;
wire \mem[4][57]~q ;
wire \mem~30_combout ;
wire \mem[3][57]~q ;
wire \mem~23_combout ;
wire \mem[2][57]~q ;
wire \mem~16_combout ;
wire \mem[1][57]~q ;
wire \mem~9_combout ;


dffeas \mem_used[7] (
	.clk(clk),
	.d(\mem_used[7]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_7),
	.prn(vcc));
defparam \mem_used[7] .is_wysiwyg = "true";
defparam \mem_used[7] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][87] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_87_0),
	.prn(vcc));
defparam \mem[0][87] .is_wysiwyg = "true";
defparam \mem[0][87] .power_up = "low";

dffeas \mem[0][88] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_88_0),
	.prn(vcc));
defparam \mem[0][88] .is_wysiwyg = "true";
defparam \mem[0][88] .power_up = "low";

dffeas \mem[0][54] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_54_0),
	.prn(vcc));
defparam \mem[0][54] .is_wysiwyg = "true";
defparam \mem[0][54] .power_up = "low";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_19_0),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][48] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_48_0),
	.prn(vcc));
defparam \mem[0][48] .is_wysiwyg = "true";
defparam \mem[0][48] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(src_data_66),
	.datab(WideOr1),
	.datac(mem_used_7),
	.datad(cp_ready),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hEFFF;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used~6 (
	.dataa(mem_used_0),
	.datab(\mem_used[2]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~6_combout ),
	.cout());
defparam \mem_used~6 .lut_mask = 16'hAACC;
defparam \mem_used~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[6]~4 (
	.dataa(src_data_66),
	.datab(mem_used_7),
	.datac(cp_ready),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[6]~4_combout ),
	.cout());
defparam \mem_used[6]~4 .lut_mask = 16'hFDFD;
defparam \mem_used[6]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[6]~5 (
	.dataa(comb),
	.datab(WideOr1),
	.datac(\mem_used[6]~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[6]~5_combout ),
	.cout());
defparam \mem_used[6]~5 .lut_mask = 16'h9696;
defparam \mem_used[6]~5 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~5_combout ),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used~8 (
	.dataa(\mem_used[1]~q ),
	.datab(\mem_used[3]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~8_combout ),
	.cout());
defparam \mem_used~8 .lut_mask = 16'hAACC;
defparam \mem_used~8 .sum_lutc_input = "datac";

dffeas \mem_used[2] (
	.clk(clk),
	.d(\mem_used~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~5_combout ),
	.q(\mem_used[2]~q ),
	.prn(vcc));
defparam \mem_used[2] .is_wysiwyg = "true";
defparam \mem_used[2] .power_up = "low";

cycloneive_lcell_comb \mem_used~10 (
	.dataa(\mem_used[2]~q ),
	.datab(\mem_used[4]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~10_combout ),
	.cout());
defparam \mem_used~10 .lut_mask = 16'hAACC;
defparam \mem_used~10 .sum_lutc_input = "datac";

dffeas \mem_used[3] (
	.clk(clk),
	.d(\mem_used~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~5_combout ),
	.q(\mem_used[3]~q ),
	.prn(vcc));
defparam \mem_used[3] .is_wysiwyg = "true";
defparam \mem_used[3] .power_up = "low";

cycloneive_lcell_comb \mem_used~9 (
	.dataa(\mem_used[3]~q ),
	.datab(\mem_used[5]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~9_combout ),
	.cout());
defparam \mem_used~9 .lut_mask = 16'hAACC;
defparam \mem_used~9 .sum_lutc_input = "datac";

dffeas \mem_used[4] (
	.clk(clk),
	.d(\mem_used~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~5_combout ),
	.q(\mem_used[4]~q ),
	.prn(vcc));
defparam \mem_used[4] .is_wysiwyg = "true";
defparam \mem_used[4] .power_up = "low";

cycloneive_lcell_comb \mem_used~7 (
	.dataa(\mem_used[4]~q ),
	.datab(\mem_used[6]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~7_combout ),
	.cout());
defparam \mem_used~7 .lut_mask = 16'hAACC;
defparam \mem_used~7 .sum_lutc_input = "datac";

dffeas \mem_used[5] (
	.clk(clk),
	.d(\mem_used~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~5_combout ),
	.q(\mem_used[5]~q ),
	.prn(vcc));
defparam \mem_used[5] .is_wysiwyg = "true";
defparam \mem_used[5] .power_up = "low";

cycloneive_lcell_comb \mem_used~3 (
	.dataa(mem_used_7),
	.datab(\write~0_combout ),
	.datac(\mem_used[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used~3_combout ),
	.cout());
defparam \mem_used~3 .lut_mask = 16'hFEFE;
defparam \mem_used~3 .sum_lutc_input = "datac";

dffeas \mem_used[6] (
	.clk(clk),
	.d(\mem_used~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~5_combout ),
	.q(\mem_used[6]~q ),
	.prn(vcc));
defparam \mem_used[6] .is_wysiwyg = "true";
defparam \mem_used[6] .power_up = "low";

cycloneive_lcell_comb \mem_used[7]~0 (
	.dataa(\mem_used[6]~q ),
	.datab(mem_used_7),
	.datac(comb),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used[7]~0_combout ),
	.cout());
defparam \mem_used[7]~0 .lut_mask = 16'hEFFE;
defparam \mem_used[7]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~1 (
	.dataa(mem_used_0),
	.datab(\mem_used[1]~q ),
	.datac(mem_87_0),
	.datad(out_valid),
	.cin(gnd),
	.combout(\mem_used[0]~1_combout ),
	.cout());
defparam \mem_used[0]~1 .lut_mask = 16'hEFFF;
defparam \mem_used[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(\write~0_combout ),
	.datab(\mem_used[0]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hEEEE;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem[7][87] (
	.clk(clk),
	.d(\mem~41_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][87]~q ),
	.prn(vcc));
defparam \mem[7][87] .is_wysiwyg = "true";
defparam \mem[7][87] .power_up = "low";

cycloneive_lcell_comb \mem~41 (
	.dataa(\mem[7][87]~q ),
	.datab(rf_source_data_87),
	.datac(gnd),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~41_combout ),
	.cout());
defparam \mem~41 .lut_mask = 16'hAACC;
defparam \mem~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always6~0 (
	.dataa(mem_used_0),
	.datab(mem_87_0),
	.datac(out_valid),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\always6~0_combout ),
	.cout());
defparam \always6~0 .lut_mask = 16'hFEFF;
defparam \always6~0 .sum_lutc_input = "datac";

dffeas \mem[6][87] (
	.clk(clk),
	.d(\mem~41_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][87]~q ),
	.prn(vcc));
defparam \mem[6][87] .is_wysiwyg = "true";
defparam \mem[6][87] .power_up = "low";

cycloneive_lcell_comb \mem~34 (
	.dataa(\mem[6][87]~q ),
	.datab(rf_source_data_87),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~34_combout ),
	.cout());
defparam \mem~34 .lut_mask = 16'hAACC;
defparam \mem~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always5~0 (
	.dataa(mem_used_0),
	.datab(mem_87_0),
	.datac(out_valid),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'hFEFF;
defparam \always5~0 .sum_lutc_input = "datac";

dffeas \mem[5][87] (
	.clk(clk),
	.d(\mem~34_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][87]~q ),
	.prn(vcc));
defparam \mem[5][87] .is_wysiwyg = "true";
defparam \mem[5][87] .power_up = "low";

cycloneive_lcell_comb \mem~27 (
	.dataa(\mem[5][87]~q ),
	.datab(rf_source_data_87),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~27_combout ),
	.cout());
defparam \mem~27 .lut_mask = 16'hAACC;
defparam \mem~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always4~0 (
	.dataa(mem_used_0),
	.datab(mem_87_0),
	.datac(out_valid),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'hFEFF;
defparam \always4~0 .sum_lutc_input = "datac";

dffeas \mem[4][87] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][87]~q ),
	.prn(vcc));
defparam \mem[4][87] .is_wysiwyg = "true";
defparam \mem[4][87] .power_up = "low";

cycloneive_lcell_comb \mem~20 (
	.dataa(\mem[4][87]~q ),
	.datab(rf_source_data_87),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~20_combout ),
	.cout());
defparam \mem~20 .lut_mask = 16'hAACC;
defparam \mem~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always3~0 (
	.dataa(mem_used_0),
	.datab(mem_87_0),
	.datac(out_valid),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\always3~0_combout ),
	.cout());
defparam \always3~0 .lut_mask = 16'hFEFF;
defparam \always3~0 .sum_lutc_input = "datac";

dffeas \mem[3][87] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][87]~q ),
	.prn(vcc));
defparam \mem[3][87] .is_wysiwyg = "true";
defparam \mem[3][87] .power_up = "low";

cycloneive_lcell_comb \mem~13 (
	.dataa(\mem[3][87]~q ),
	.datab(rf_source_data_87),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~13_combout ),
	.cout());
defparam \mem~13 .lut_mask = 16'hAACC;
defparam \mem~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(mem_used_0),
	.datab(mem_87_0),
	.datac(out_valid),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hFEFF;
defparam \always2~0 .sum_lutc_input = "datac";

dffeas \mem[2][87] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][87]~q ),
	.prn(vcc));
defparam \mem[2][87] .is_wysiwyg = "true";
defparam \mem[2][87] .power_up = "low";

cycloneive_lcell_comb \mem~6 (
	.dataa(\mem[2][87]~q ),
	.datab(rf_source_data_87),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~6_combout ),
	.cout());
defparam \mem~6 .lut_mask = 16'hAACC;
defparam \mem~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(mem_used_0),
	.datab(mem_87_0),
	.datac(out_valid),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hFEFF;
defparam \always1~0 .sum_lutc_input = "datac";

dffeas \mem[1][87] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][87]~q ),
	.prn(vcc));
defparam \mem[1][87] .is_wysiwyg = "true";
defparam \mem[1][87] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][87]~q ),
	.datab(rf_source_data_87),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(mem_87_0),
	.datab(out_valid),
	.datac(gnd),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hEEFF;
defparam \always0~0 .sum_lutc_input = "datac";

dffeas \mem[7][88] (
	.clk(clk),
	.d(\mem~42_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][88]~q ),
	.prn(vcc));
defparam \mem[7][88] .is_wysiwyg = "true";
defparam \mem[7][88] .power_up = "low";

cycloneive_lcell_comb \mem~42 (
	.dataa(\mem[7][88]~q ),
	.datab(out_endofpacket),
	.datac(gnd),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~42_combout ),
	.cout());
defparam \mem~42 .lut_mask = 16'hAACC;
defparam \mem~42 .sum_lutc_input = "datac";

dffeas \mem[6][88] (
	.clk(clk),
	.d(\mem~42_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][88]~q ),
	.prn(vcc));
defparam \mem[6][88] .is_wysiwyg = "true";
defparam \mem[6][88] .power_up = "low";

cycloneive_lcell_comb \mem~35 (
	.dataa(\mem[6][88]~q ),
	.datab(out_endofpacket),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~35_combout ),
	.cout());
defparam \mem~35 .lut_mask = 16'hAACC;
defparam \mem~35 .sum_lutc_input = "datac";

dffeas \mem[5][88] (
	.clk(clk),
	.d(\mem~35_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][88]~q ),
	.prn(vcc));
defparam \mem[5][88] .is_wysiwyg = "true";
defparam \mem[5][88] .power_up = "low";

cycloneive_lcell_comb \mem~28 (
	.dataa(\mem[5][88]~q ),
	.datab(out_endofpacket),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~28_combout ),
	.cout());
defparam \mem~28 .lut_mask = 16'hAACC;
defparam \mem~28 .sum_lutc_input = "datac";

dffeas \mem[4][88] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][88]~q ),
	.prn(vcc));
defparam \mem[4][88] .is_wysiwyg = "true";
defparam \mem[4][88] .power_up = "low";

cycloneive_lcell_comb \mem~21 (
	.dataa(\mem[4][88]~q ),
	.datab(out_endofpacket),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~21_combout ),
	.cout());
defparam \mem~21 .lut_mask = 16'hAACC;
defparam \mem~21 .sum_lutc_input = "datac";

dffeas \mem[3][88] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][88]~q ),
	.prn(vcc));
defparam \mem[3][88] .is_wysiwyg = "true";
defparam \mem[3][88] .power_up = "low";

cycloneive_lcell_comb \mem~14 (
	.dataa(\mem[3][88]~q ),
	.datab(out_endofpacket),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~14_combout ),
	.cout());
defparam \mem~14 .lut_mask = 16'hAACC;
defparam \mem~14 .sum_lutc_input = "datac";

dffeas \mem[2][88] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][88]~q ),
	.prn(vcc));
defparam \mem[2][88] .is_wysiwyg = "true";
defparam \mem[2][88] .power_up = "low";

cycloneive_lcell_comb \mem~7 (
	.dataa(\mem[2][88]~q ),
	.datab(out_endofpacket),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~7_combout ),
	.cout());
defparam \mem~7 .lut_mask = 16'hAACC;
defparam \mem~7 .sum_lutc_input = "datac";

dffeas \mem[1][88] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][88]~q ),
	.prn(vcc));
defparam \mem[1][88] .is_wysiwyg = "true";
defparam \mem[1][88] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][88]~q ),
	.datab(out_endofpacket),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[7][85] (
	.clk(clk),
	.d(\mem~43_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][85]~q ),
	.prn(vcc));
defparam \mem[7][85] .is_wysiwyg = "true";
defparam \mem[7][85] .power_up = "low";

cycloneive_lcell_comb \mem~43 (
	.dataa(\mem[7][85]~q ),
	.datab(saved_grant_0),
	.datac(saved_grant_1),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~43_combout ),
	.cout());
defparam \mem~43 .lut_mask = 16'hFAFC;
defparam \mem~43 .sum_lutc_input = "datac";

dffeas \mem[6][54] (
	.clk(clk),
	.d(\mem~43_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][54]~q ),
	.prn(vcc));
defparam \mem[6][54] .is_wysiwyg = "true";
defparam \mem[6][54] .power_up = "low";

cycloneive_lcell_comb \mem~36 (
	.dataa(\mem[6][54]~q ),
	.datab(saved_grant_0),
	.datac(saved_grant_1),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~36_combout ),
	.cout());
defparam \mem~36 .lut_mask = 16'hFAFC;
defparam \mem~36 .sum_lutc_input = "datac";

dffeas \mem[5][54] (
	.clk(clk),
	.d(\mem~36_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][54]~q ),
	.prn(vcc));
defparam \mem[5][54] .is_wysiwyg = "true";
defparam \mem[5][54] .power_up = "low";

cycloneive_lcell_comb \mem~29 (
	.dataa(\mem[5][54]~q ),
	.datab(saved_grant_0),
	.datac(saved_grant_1),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~29_combout ),
	.cout());
defparam \mem~29 .lut_mask = 16'hFAFC;
defparam \mem~29 .sum_lutc_input = "datac";

dffeas \mem[4][54] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][54]~q ),
	.prn(vcc));
defparam \mem[4][54] .is_wysiwyg = "true";
defparam \mem[4][54] .power_up = "low";

cycloneive_lcell_comb \mem~22 (
	.dataa(\mem[4][54]~q ),
	.datab(saved_grant_0),
	.datac(saved_grant_1),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~22_combout ),
	.cout());
defparam \mem~22 .lut_mask = 16'hFAFC;
defparam \mem~22 .sum_lutc_input = "datac";

dffeas \mem[3][54] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][54]~q ),
	.prn(vcc));
defparam \mem[3][54] .is_wysiwyg = "true";
defparam \mem[3][54] .power_up = "low";

cycloneive_lcell_comb \mem~15 (
	.dataa(\mem[3][54]~q ),
	.datab(saved_grant_0),
	.datac(saved_grant_1),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~15_combout ),
	.cout());
defparam \mem~15 .lut_mask = 16'hFAFC;
defparam \mem~15 .sum_lutc_input = "datac";

dffeas \mem[2][54] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][54]~q ),
	.prn(vcc));
defparam \mem[2][54] .is_wysiwyg = "true";
defparam \mem[2][54] .power_up = "low";

cycloneive_lcell_comb \mem~8 (
	.dataa(\mem[2][54]~q ),
	.datab(saved_grant_0),
	.datac(saved_grant_1),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~8_combout ),
	.cout());
defparam \mem~8 .lut_mask = 16'hFAFC;
defparam \mem~8 .sum_lutc_input = "datac";

dffeas \mem[1][54] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][54]~q ),
	.prn(vcc));
defparam \mem[1][54] .is_wysiwyg = "true";
defparam \mem[1][54] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][54]~q ),
	.datab(saved_grant_0),
	.datac(saved_grant_1),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hFAFC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[7][19] (
	.clk(clk),
	.d(\mem~45_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][19]~q ),
	.prn(vcc));
defparam \mem[7][19] .is_wysiwyg = "true";
defparam \mem[7][19] .power_up = "low";

cycloneive_lcell_comb \mem~45 (
	.dataa(\mem[7][19]~q ),
	.datab(use_reg),
	.datac(address_reg_1),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~45_combout ),
	.cout());
defparam \mem~45 .lut_mask = 16'hFAFC;
defparam \mem~45 .sum_lutc_input = "datac";

dffeas \mem[6][19] (
	.clk(clk),
	.d(\mem~45_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][19]~q ),
	.prn(vcc));
defparam \mem[6][19] .is_wysiwyg = "true";
defparam \mem[6][19] .power_up = "low";

cycloneive_lcell_comb \mem~38 (
	.dataa(\mem[6][19]~q ),
	.datab(use_reg),
	.datac(address_reg_1),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~38_combout ),
	.cout());
defparam \mem~38 .lut_mask = 16'hFAFC;
defparam \mem~38 .sum_lutc_input = "datac";

dffeas \mem[5][19] (
	.clk(clk),
	.d(\mem~38_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][19]~q ),
	.prn(vcc));
defparam \mem[5][19] .is_wysiwyg = "true";
defparam \mem[5][19] .power_up = "low";

cycloneive_lcell_comb \mem~31 (
	.dataa(\mem[5][19]~q ),
	.datab(use_reg),
	.datac(address_reg_1),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~31_combout ),
	.cout());
defparam \mem~31 .lut_mask = 16'hFAFC;
defparam \mem~31 .sum_lutc_input = "datac";

dffeas \mem[4][19] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][19]~q ),
	.prn(vcc));
defparam \mem[4][19] .is_wysiwyg = "true";
defparam \mem[4][19] .power_up = "low";

cycloneive_lcell_comb \mem~24 (
	.dataa(\mem[4][19]~q ),
	.datab(use_reg),
	.datac(address_reg_1),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~24_combout ),
	.cout());
defparam \mem~24 .lut_mask = 16'hFAFC;
defparam \mem~24 .sum_lutc_input = "datac";

dffeas \mem[3][19] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][19]~q ),
	.prn(vcc));
defparam \mem[3][19] .is_wysiwyg = "true";
defparam \mem[3][19] .power_up = "low";

cycloneive_lcell_comb \mem~17 (
	.dataa(\mem[3][19]~q ),
	.datab(use_reg),
	.datac(address_reg_1),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~17_combout ),
	.cout());
defparam \mem~17 .lut_mask = 16'hFAFC;
defparam \mem~17 .sum_lutc_input = "datac";

dffeas \mem[2][19] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][19]~q ),
	.prn(vcc));
defparam \mem[2][19] .is_wysiwyg = "true";
defparam \mem[2][19] .power_up = "low";

cycloneive_lcell_comb \mem~10 (
	.dataa(\mem[2][19]~q ),
	.datab(use_reg),
	.datac(address_reg_1),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~10_combout ),
	.cout());
defparam \mem~10 .lut_mask = 16'hFAFC;
defparam \mem~10 .sum_lutc_input = "datac";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][19]~q ),
	.datab(use_reg),
	.datac(address_reg_1),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hFAFC;
defparam \mem~3 .sum_lutc_input = "datac";

dffeas \mem[7][66] (
	.clk(clk),
	.d(\mem~46_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][66]~q ),
	.prn(vcc));
defparam \mem[7][66] .is_wysiwyg = "true";
defparam \mem[7][66] .power_up = "low";

cycloneive_lcell_comb \mem~46 (
	.dataa(\mem[7][66]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~46_combout ),
	.cout());
defparam \mem~46 .lut_mask = 16'hAACC;
defparam \mem~46 .sum_lutc_input = "datac";

dffeas \mem[6][66] (
	.clk(clk),
	.d(\mem~46_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][66]~q ),
	.prn(vcc));
defparam \mem[6][66] .is_wysiwyg = "true";
defparam \mem[6][66] .power_up = "low";

cycloneive_lcell_comb \mem~39 (
	.dataa(\mem[6][66]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~39_combout ),
	.cout());
defparam \mem~39 .lut_mask = 16'hAACC;
defparam \mem~39 .sum_lutc_input = "datac";

dffeas \mem[5][66] (
	.clk(clk),
	.d(\mem~39_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][66]~q ),
	.prn(vcc));
defparam \mem[5][66] .is_wysiwyg = "true";
defparam \mem[5][66] .power_up = "low";

cycloneive_lcell_comb \mem~32 (
	.dataa(\mem[5][66]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~32_combout ),
	.cout());
defparam \mem~32 .lut_mask = 16'hAACC;
defparam \mem~32 .sum_lutc_input = "datac";

dffeas \mem[4][66] (
	.clk(clk),
	.d(\mem~32_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][66]~q ),
	.prn(vcc));
defparam \mem[4][66] .is_wysiwyg = "true";
defparam \mem[4][66] .power_up = "low";

cycloneive_lcell_comb \mem~25 (
	.dataa(\mem[4][66]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~25_combout ),
	.cout());
defparam \mem~25 .lut_mask = 16'hAACC;
defparam \mem~25 .sum_lutc_input = "datac";

dffeas \mem[3][66] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][66]~q ),
	.prn(vcc));
defparam \mem[3][66] .is_wysiwyg = "true";
defparam \mem[3][66] .power_up = "low";

cycloneive_lcell_comb \mem~18 (
	.dataa(\mem[3][66]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~18_combout ),
	.cout());
defparam \mem~18 .lut_mask = 16'hAACC;
defparam \mem~18 .sum_lutc_input = "datac";

dffeas \mem[2][66] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][66]~q ),
	.prn(vcc));
defparam \mem[2][66] .is_wysiwyg = "true";
defparam \mem[2][66] .power_up = "low";

cycloneive_lcell_comb \mem~11 (
	.dataa(\mem[2][66]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~11_combout ),
	.cout());
defparam \mem~11 .lut_mask = 16'hAACC;
defparam \mem~11 .sum_lutc_input = "datac";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[1][66]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hAACC;
defparam \mem~4 .sum_lutc_input = "datac";

dffeas \mem[7][48] (
	.clk(clk),
	.d(\mem~47_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][48]~q ),
	.prn(vcc));
defparam \mem[7][48] .is_wysiwyg = "true";
defparam \mem[7][48] .power_up = "low";

cycloneive_lcell_comb \mem~47 (
	.dataa(\mem[7][48]~q ),
	.datab(src_data_66),
	.datac(gnd),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~47_combout ),
	.cout());
defparam \mem~47 .lut_mask = 16'hAACC;
defparam \mem~47 .sum_lutc_input = "datac";

dffeas \mem[6][48] (
	.clk(clk),
	.d(\mem~47_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][48]~q ),
	.prn(vcc));
defparam \mem[6][48] .is_wysiwyg = "true";
defparam \mem[6][48] .power_up = "low";

cycloneive_lcell_comb \mem~40 (
	.dataa(\mem[6][48]~q ),
	.datab(src_data_66),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~40_combout ),
	.cout());
defparam \mem~40 .lut_mask = 16'hAACC;
defparam \mem~40 .sum_lutc_input = "datac";

dffeas \mem[5][48] (
	.clk(clk),
	.d(\mem~40_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][48]~q ),
	.prn(vcc));
defparam \mem[5][48] .is_wysiwyg = "true";
defparam \mem[5][48] .power_up = "low";

cycloneive_lcell_comb \mem~33 (
	.dataa(\mem[5][48]~q ),
	.datab(src_data_66),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~33_combout ),
	.cout());
defparam \mem~33 .lut_mask = 16'hAACC;
defparam \mem~33 .sum_lutc_input = "datac";

dffeas \mem[4][48] (
	.clk(clk),
	.d(\mem~33_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][48]~q ),
	.prn(vcc));
defparam \mem[4][48] .is_wysiwyg = "true";
defparam \mem[4][48] .power_up = "low";

cycloneive_lcell_comb \mem~26 (
	.dataa(\mem[4][48]~q ),
	.datab(src_data_66),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~26_combout ),
	.cout());
defparam \mem~26 .lut_mask = 16'hAACC;
defparam \mem~26 .sum_lutc_input = "datac";

dffeas \mem[3][48] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][48]~q ),
	.prn(vcc));
defparam \mem[3][48] .is_wysiwyg = "true";
defparam \mem[3][48] .power_up = "low";

cycloneive_lcell_comb \mem~19 (
	.dataa(\mem[3][48]~q ),
	.datab(src_data_66),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~19_combout ),
	.cout());
defparam \mem~19 .lut_mask = 16'hAACC;
defparam \mem~19 .sum_lutc_input = "datac";

dffeas \mem[2][48] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][48]~q ),
	.prn(vcc));
defparam \mem[2][48] .is_wysiwyg = "true";
defparam \mem[2][48] .power_up = "low";

cycloneive_lcell_comb \mem~12 (
	.dataa(\mem[2][48]~q ),
	.datab(src_data_66),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~12_combout ),
	.cout());
defparam \mem~12 .lut_mask = 16'hAACC;
defparam \mem~12 .sum_lutc_input = "datac";

dffeas \mem[1][48] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][48]~q ),
	.prn(vcc));
defparam \mem[1][48] .is_wysiwyg = "true";
defparam \mem[1][48] .power_up = "low";

cycloneive_lcell_comb \mem~5 (
	.dataa(\mem[1][48]~q ),
	.datab(src_data_66),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~5_combout ),
	.cout());
defparam \mem~5 .lut_mask = 16'hAACC;
defparam \mem~5 .sum_lutc_input = "datac";

dffeas \mem[7][57] (
	.clk(clk),
	.d(\mem~48_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][57]~q ),
	.prn(vcc));
defparam \mem[7][57] .is_wysiwyg = "true";
defparam \mem[7][57] .power_up = "low";

cycloneive_lcell_comb \mem~48 (
	.dataa(\mem[7][57]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~48_combout ),
	.cout());
defparam \mem~48 .lut_mask = 16'hAAFF;
defparam \mem~48 .sum_lutc_input = "datac";

dffeas \mem[6][57] (
	.clk(clk),
	.d(\mem~48_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][57]~q ),
	.prn(vcc));
defparam \mem[6][57] .is_wysiwyg = "true";
defparam \mem[6][57] .power_up = "low";

cycloneive_lcell_comb \mem~44 (
	.dataa(\mem[6][57]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~44_combout ),
	.cout());
defparam \mem~44 .lut_mask = 16'hAAFF;
defparam \mem~44 .sum_lutc_input = "datac";

dffeas \mem[5][57] (
	.clk(clk),
	.d(\mem~44_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][57]~q ),
	.prn(vcc));
defparam \mem[5][57] .is_wysiwyg = "true";
defparam \mem[5][57] .power_up = "low";

cycloneive_lcell_comb \mem~37 (
	.dataa(\mem[5][57]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~37_combout ),
	.cout());
defparam \mem~37 .lut_mask = 16'hAAFF;
defparam \mem~37 .sum_lutc_input = "datac";

dffeas \mem[4][57] (
	.clk(clk),
	.d(\mem~37_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][57]~q ),
	.prn(vcc));
defparam \mem[4][57] .is_wysiwyg = "true";
defparam \mem[4][57] .power_up = "low";

cycloneive_lcell_comb \mem~30 (
	.dataa(\mem[4][57]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~30_combout ),
	.cout());
defparam \mem~30 .lut_mask = 16'hAAFF;
defparam \mem~30 .sum_lutc_input = "datac";

dffeas \mem[3][57] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][57]~q ),
	.prn(vcc));
defparam \mem[3][57] .is_wysiwyg = "true";
defparam \mem[3][57] .power_up = "low";

cycloneive_lcell_comb \mem~23 (
	.dataa(\mem[3][57]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~23_combout ),
	.cout());
defparam \mem~23 .lut_mask = 16'hAAFF;
defparam \mem~23 .sum_lutc_input = "datac";

dffeas \mem[2][57] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][57]~q ),
	.prn(vcc));
defparam \mem[2][57] .is_wysiwyg = "true";
defparam \mem[2][57] .power_up = "low";

cycloneive_lcell_comb \mem~16 (
	.dataa(\mem[2][57]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~16_combout ),
	.cout());
defparam \mem~16 .lut_mask = 16'hAAFF;
defparam \mem~16 .sum_lutc_input = "datac";

dffeas \mem[1][57] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][57]~q ),
	.prn(vcc));
defparam \mem[1][57] .is_wysiwyg = "true";
defparam \mem[1][57] .power_up = "low";

cycloneive_lcell_comb \mem~9 (
	.dataa(\mem[1][57]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~9_combout ),
	.cout());
defparam \mem~9 .lut_mask = 16'hAAFF;
defparam \mem~9 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_14 (
	clk,
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~1 (
	.dataa(sink_ready),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~1_combout ),
	.cout());
defparam \mem_used[0]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~1 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(mem_used_1),
	.datab(sink_ready1),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hACFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_15 (
	reset,
	mem_used_0,
	mem_105_0,
	read_latency_shift_reg_0,
	mem_used_01,
	rp_valid,
	in_ready,
	av_readdata_pre_0,
	out_data_0,
	av_readdata_pre_1,
	out_data_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	mem_used_0;
input 	mem_105_0;
input 	read_latency_shift_reg_0;
output 	mem_used_01;
input 	rp_valid;
input 	in_ready;
input 	av_readdata_pre_0;
output 	out_data_0;
input 	av_readdata_pre_1;
output 	out_data_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[0][0]~q ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[0][1]~q ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_01),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \out_data[0]~0 (
	.dataa(\mem[0][0]~q ),
	.datab(av_readdata_pre_0),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_0),
	.cout());
defparam \out_data[0]~0 .lut_mask = 16'hEFFE;
defparam \out_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[1]~1 (
	.dataa(\mem[0][1]~q ),
	.datab(av_readdata_pre_1),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_1),
	.cout());
defparam \out_data[1]~1 .lut_mask = 16'hEFFE;
defparam \out_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(mem_used_0),
	.datab(mem_105_0),
	.datac(in_ready),
	.datad(rp_valid),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h7FFF;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[1]~q ),
	.datab(read_latency_shift_reg_0),
	.datac(mem_used_01),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~0 (
	.dataa(\mem_used[1]~q ),
	.datab(mem_used_01),
	.datac(read_latency_shift_reg_0),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~0_combout ),
	.cout());
defparam \mem_used[0]~0 .lut_mask = 16'hFDFE;
defparam \mem_used[0]~0 .sum_lutc_input = "datac";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][0]~q ),
	.datab(av_readdata_pre_0),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hAAFF;
defparam \always0~0 .sum_lutc_input = "datac";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][0]~q ),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][1]~q ),
	.datab(av_readdata_pre_1),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][1]~q ),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

endmodule

module niosII_altera_avalon_sc_fifo_16 (
	out_data_toggle_flopped,
	dreg_0,
	mem_used_1,
	wire_pfdena_reg_ena,
	out_data_buffer_65,
	reset,
	rst1,
	mem_used_0,
	out_data_buffer_66,
	out_data_buffer_105,
	out_data_buffer_64,
	mem_105_0,
	sink_ready,
	clk)/* synthesis synthesis_greybox=1 */;
input 	out_data_toggle_flopped;
input 	dreg_0;
output 	mem_used_1;
input 	wire_pfdena_reg_ena;
input 	out_data_buffer_65;
input 	reset;
input 	rst1;
output 	mem_used_0;
input 	out_data_buffer_66;
input 	out_data_buffer_105;
input 	out_data_buffer_64;
output 	mem_105_0;
input 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem[1][105]~q ;
wire \mem~1_combout ;
wire \mem[0][105]~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem[0][105]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(out_data_buffer_65),
	.datab(out_data_buffer_105),
	.datac(gnd),
	.datad(out_data_buffer_64),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hEEFF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(mem_used_0),
	.datab(out_data_buffer_66),
	.datac(\mem~0_combout ),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(rst1),
	.datab(\mem_used[1]~0_combout ),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hEFFE;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(mem_used_1),
	.datac(mem_used_0),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(wire_pfdena_reg_ena),
	.datab(rst1),
	.datac(out_data_buffer_66),
	.datad(\mem~0_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(mem_used_0),
	.datac(mem_used_1),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(mem_used_1),
	.datab(wire_pfdena_reg_ena),
	.datac(\mem~0_combout ),
	.datad(\mem[1][105]~q ),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hFFFE;
defparam \mem~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][105]~2 (
	.dataa(\mem~1_combout ),
	.datab(mem_105_0),
	.datac(mem_used_0),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\mem[0][105]~2_combout ),
	.cout());
defparam \mem[0][105]~2 .lut_mask = 16'hEFFE;
defparam \mem[0][105]~2 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_sc_fifo_17 (
	clk,
	reset,
	uav_read,
	hold_waitrequest,
	Equal4,
	read_latency_shift_reg_0,
	mem_used_1,
	wait_latency_counter_1,
	av_waitrequest_generated,
	period_l_wr_strobe)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	uav_read;
input 	hold_waitrequest;
input 	Equal4;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	wait_latency_counter_1;
input 	av_waitrequest_generated;
input 	period_l_wr_strobe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(uav_read),
	.datac(av_waitrequest_generated),
	.datad(period_l_wr_strobe),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(hold_waitrequest),
	.datab(uav_read),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(Equal4),
	.datab(av_waitrequest_generated),
	.datac(\mem_used[1]~0_combout ),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module niosII_altera_avalon_st_handshake_clock_crosser (
	wire_pll7_clk_0,
	W_alu_result_2,
	r_sync_rst,
	uav_read,
	cp_valid,
	d_writedata_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	altera_reset_synchronizer_int_chain_out,
	Equal13,
	in_data_toggle,
	dreg_0,
	d_writedata_10,
	uav_write,
	out_data_toggle_flopped,
	dreg_01,
	av_waitrequest,
	mem_used_1,
	out_data_buffer_66,
	out_data_buffer_38,
	out_data_buffer_7,
	out_data_buffer_65,
	out_data_buffer_105,
	out_data_buffer_64,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_10,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_2;
input 	r_sync_rst;
input 	uav_read;
input 	cp_valid;
input 	d_writedata_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal13;
output 	in_data_toggle;
output 	dreg_0;
input 	d_writedata_10;
input 	uav_write;
output 	out_data_toggle_flopped;
output 	dreg_01;
input 	av_waitrequest;
input 	mem_used_1;
output 	out_data_buffer_66;
output 	out_data_buffer_38;
output 	out_data_buffer_7;
output 	out_data_buffer_65;
output 	out_data_buffer_105;
output 	out_data_buffer_64;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_10;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_avalon_st_clock_crosser_7 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,uav_read,uav_write,uav_write,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,W_alu_result_2,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_10,gnd,gnd,d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.in_reset(r_sync_rst),
	.cp_valid(cp_valid),
	.out_reset(altera_reset_synchronizer_int_chain_out),
	.Equal13(Equal13),
	.in_data_toggle1(in_data_toggle),
	.dreg_0(dreg_0),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_01(dreg_01),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_1),
	.out_data_buffer_66(out_data_buffer_66),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_65(out_data_buffer_65),
	.out_data_buffer_105(out_data_buffer_105),
	.out_data_buffer_64(out_data_buffer_64),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_6(out_data_buffer_6),
	.clk_clk(clk_clk));

endmodule

module niosII_altera_avalon_st_handshake_clock_crosser_1 (
	wire_pll7_clk_0,
	W_alu_result_6,
	W_alu_result_10,
	W_alu_result_5,
	W_alu_result_7,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	r_sync_rst,
	r_sync_rst1,
	saved_grant_0,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_10,
	uav_read,
	out_data_buffer_0,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	last_cycle,
	out_data_buffer_105,
	out_data_buffer_46,
	out_data_buffer_65,
	out_data_buffer_7,
	d_writedata_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	Equal1,
	src12_valid,
	in_ready,
	out_data_buffer_66,
	out_data_buffer_64,
	d_writedata_10,
	out_data_buffer_6,
	d_writedata_8,
	d_writedata_9,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	uav_write,
	out_data_buffer_5,
	out_data_buffer_4,
	out_data_buffer_3,
	out_data_buffer_2,
	out_data_buffer_1,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_12,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_9,
	out_data_buffer_8)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_6;
input 	W_alu_result_10;
input 	W_alu_result_5;
input 	W_alu_result_7;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	r_sync_rst;
input 	r_sync_rst1;
input 	saved_grant_0;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_10;
input 	uav_read;
output 	out_data_buffer_0;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	out_valid;
input 	last_cycle;
output 	out_data_buffer_105;
output 	out_data_buffer_46;
output 	out_data_buffer_65;
output 	out_data_buffer_7;
input 	d_writedata_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	Equal1;
input 	src12_valid;
output 	in_ready;
output 	out_data_buffer_66;
output 	out_data_buffer_64;
input 	d_writedata_10;
output 	out_data_buffer_6;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	uav_write;
output 	out_data_buffer_5;
output 	out_data_buffer_4;
output 	out_data_buffer_3;
output 	out_data_buffer_2;
output 	out_data_buffer_1;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_12;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_9;
output 	out_data_buffer_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_avalon_st_clock_crosser clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,uav_read,uav_write,uav_write,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,W_alu_result_10,
W_alu_result_9,W_alu_result_8,W_alu_result_7,W_alu_result_6,W_alu_result_5,W_alu_result_4,W_alu_result_3,W_alu_result_2,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_15,d_writedata_14,d_writedata_13,d_writedata_12,d_writedata_11,
d_writedata_10,d_writedata_9,d_writedata_8,d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.in_reset(r_sync_rst),
	.out_reset(r_sync_rst1),
	.saved_grant_0(saved_grant_0),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(out_data_buffer_39),
	.out_data_buffer_40(out_data_buffer_40),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid),
	.last_cycle(last_cycle),
	.out_data_buffer_105(out_data_buffer_105),
	.out_data_buffer_46(out_data_buffer_46),
	.out_data_buffer_65(out_data_buffer_65),
	.out_data_buffer_7(out_data_buffer_7),
	.Equal1(Equal1),
	.src12_valid(src12_valid),
	.in_ready(in_ready),
	.out_data_buffer_66(out_data_buffer_66),
	.out_data_buffer_64(out_data_buffer_64),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_41(out_data_buffer_41),
	.out_data_buffer_42(out_data_buffer_42),
	.out_data_buffer_43(out_data_buffer_43),
	.out_data_buffer_44(out_data_buffer_44),
	.out_data_buffer_45(out_data_buffer_45),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_8(out_data_buffer_8));

endmodule

module niosII_altera_avalon_st_clock_crosser (
	wire_pll7_clk_0,
	in_data,
	in_reset,
	out_reset,
	saved_grant_0,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_10,
	out_data_buffer_0,
	out_data_toggle_flopped1,
	dreg_0,
	out_valid1,
	last_cycle,
	out_data_buffer_105,
	out_data_buffer_46,
	out_data_buffer_65,
	out_data_buffer_7,
	Equal1,
	src12_valid,
	in_ready,
	out_data_buffer_66,
	out_data_buffer_64,
	out_data_buffer_6,
	out_data_buffer_5,
	out_data_buffer_4,
	out_data_buffer_3,
	out_data_buffer_2,
	out_data_buffer_1,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_12,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_9,
	out_data_buffer_8)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	[120:0] in_data;
input 	in_reset;
input 	out_reset;
input 	saved_grant_0;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_10;
output 	out_data_buffer_0;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	out_valid1;
input 	last_cycle;
output 	out_data_buffer_105;
output 	out_data_buffer_46;
output 	out_data_buffer_65;
output 	out_data_buffer_7;
input 	Equal1;
input 	src12_valid;
output 	in_ready;
output 	out_data_buffer_66;
output 	out_data_buffer_64;
output 	out_data_buffer_6;
output 	out_data_buffer_5;
output 	out_data_buffer_4;
output 	out_data_buffer_3;
output 	out_data_buffer_2;
output 	out_data_buffer_1;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_12;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_9;
output 	out_data_buffer_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_to_in_synchronizer|dreg[0]~q ;
wire \in_data_toggle~2_combout ;
wire \in_data_toggle~q ;
wire \take_in_data~2_combout ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[39]~q ;
wire \in_data_buffer[40]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[0]~q ;
wire \out_data_toggle_flopped~0_combout ;
wire \in_data_buffer[105]~q ;
wire \in_data_buffer[46]~q ;
wire \in_data_buffer[65]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[66]~q ;
wire \in_data_buffer[64]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[41]~q ;
wire \in_data_buffer[42]~q ;
wire \in_data_buffer[43]~q ;
wire \in_data_buffer[44]~q ;
wire \in_data_buffer[45]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[8]~q ;


niosII_altera_std_synchronizer_nocut_1 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(\out_to_in_synchronizer|dreg[0]~q ));

niosII_altera_std_synchronizer_nocut in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.dreg_0(dreg_0),
	.din(\in_data_toggle~q ));

dffeas \out_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[39] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[39]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_39),
	.prn(vcc));
defparam \out_data_buffer[39] .is_wysiwyg = "true";
defparam \out_data_buffer[39] .power_up = "low";

dffeas \out_data_buffer[40] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[40]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_40),
	.prn(vcc));
defparam \out_data_buffer[40] .is_wysiwyg = "true";
defparam \out_data_buffer[40] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[105] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[105]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_105),
	.prn(vcc));
defparam \out_data_buffer[105] .is_wysiwyg = "true";
defparam \out_data_buffer[105] .power_up = "low";

dffeas \out_data_buffer[46] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[46]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_46),
	.prn(vcc));
defparam \out_data_buffer[46] .is_wysiwyg = "true";
defparam \out_data_buffer[46] .power_up = "low";

dffeas \out_data_buffer[65] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[65]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_65),
	.prn(vcc));
defparam \out_data_buffer[65] .is_wysiwyg = "true";
defparam \out_data_buffer[65] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

cycloneive_lcell_comb \in_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_data_toggle~q ),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(in_ready),
	.cout());
defparam \in_ready~0 .lut_mask = 16'h0FF0;
defparam \in_ready~0 .sum_lutc_input = "datac";

dffeas \out_data_buffer[66] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[66]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_66),
	.prn(vcc));
defparam \out_data_buffer[66] .is_wysiwyg = "true";
defparam \out_data_buffer[66] .power_up = "low";

dffeas \out_data_buffer[64] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[64]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_64),
	.prn(vcc));
defparam \out_data_buffer[64] .is_wysiwyg = "true";
defparam \out_data_buffer[64] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[41] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[41]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_41),
	.prn(vcc));
defparam \out_data_buffer[41] .is_wysiwyg = "true";
defparam \out_data_buffer[41] .power_up = "low";

dffeas \out_data_buffer[42] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[42]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_42),
	.prn(vcc));
defparam \out_data_buffer[42] .is_wysiwyg = "true";
defparam \out_data_buffer[42] .power_up = "low";

dffeas \out_data_buffer[43] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[43]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_43),
	.prn(vcc));
defparam \out_data_buffer[43] .is_wysiwyg = "true";
defparam \out_data_buffer[43] .power_up = "low";

dffeas \out_data_buffer[44] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[44]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_44),
	.prn(vcc));
defparam \out_data_buffer[44] .is_wysiwyg = "true";
defparam \out_data_buffer[44] .power_up = "low";

dffeas \out_data_buffer[45] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[45]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_45),
	.prn(vcc));
defparam \out_data_buffer[45] .is_wysiwyg = "true";
defparam \out_data_buffer[45] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~2 (
	.dataa(\in_data_toggle~q ),
	.datab(\out_to_in_synchronizer|dreg[0]~q ),
	.datac(Equal1),
	.datad(src12_valid),
	.cin(gnd),
	.combout(\in_data_toggle~2_combout ),
	.cout());
defparam \in_data_toggle~2 .lut_mask = 16'hBFFB;
defparam \in_data_toggle~2 .sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~2_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_data_toggle~q ),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb \take_in_data~2 (
	.dataa(\in_data_toggle~q ),
	.datab(\out_to_in_synchronizer|dreg[0]~q ),
	.datac(Equal1),
	.datad(src12_valid),
	.cin(gnd),
	.combout(\take_in_data~2_combout ),
	.cout());
defparam \take_in_data~2 .lut_mask = 16'hFFF6;
defparam \take_in_data~2 .sum_lutc_input = "datac";

dffeas \in_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[39] (
	.clk(wire_pll7_clk_0),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[39]~q ),
	.prn(vcc));
defparam \in_data_buffer[39] .is_wysiwyg = "true";
defparam \in_data_buffer[39] .power_up = "low";

dffeas \in_data_buffer[40] (
	.clk(wire_pll7_clk_0),
	.d(in_data[40]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[40]~q ),
	.prn(vcc));
defparam \in_data_buffer[40] .is_wysiwyg = "true";
defparam \in_data_buffer[40] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(dreg_0),
	.datab(out_data_toggle_flopped1),
	.datac(saved_grant_0),
	.datad(last_cycle),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[105] (
	.clk(wire_pll7_clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[105]~q ),
	.prn(vcc));
defparam \in_data_buffer[105] .is_wysiwyg = "true";
defparam \in_data_buffer[105] .power_up = "low";

dffeas \in_data_buffer[46] (
	.clk(wire_pll7_clk_0),
	.d(in_data[46]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[46]~q ),
	.prn(vcc));
defparam \in_data_buffer[46] .is_wysiwyg = "true";
defparam \in_data_buffer[46] .power_up = "low";

dffeas \in_data_buffer[65] (
	.clk(wire_pll7_clk_0),
	.d(in_data[65]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[65]~q ),
	.prn(vcc));
defparam \in_data_buffer[65] .is_wysiwyg = "true";
defparam \in_data_buffer[65] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[66] (
	.clk(wire_pll7_clk_0),
	.d(in_data[66]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[66]~q ),
	.prn(vcc));
defparam \in_data_buffer[66] .is_wysiwyg = "true";
defparam \in_data_buffer[66] .power_up = "low";

dffeas \in_data_buffer[64] (
	.clk(wire_pll7_clk_0),
	.d(in_data[65]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[64]~q ),
	.prn(vcc));
defparam \in_data_buffer[64] .is_wysiwyg = "true";
defparam \in_data_buffer[64] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[41] (
	.clk(wire_pll7_clk_0),
	.d(in_data[41]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[41]~q ),
	.prn(vcc));
defparam \in_data_buffer[41] .is_wysiwyg = "true";
defparam \in_data_buffer[41] .power_up = "low";

dffeas \in_data_buffer[42] (
	.clk(wire_pll7_clk_0),
	.d(in_data[42]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[42]~q ),
	.prn(vcc));
defparam \in_data_buffer[42] .is_wysiwyg = "true";
defparam \in_data_buffer[42] .power_up = "low";

dffeas \in_data_buffer[43] (
	.clk(wire_pll7_clk_0),
	.d(in_data[43]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[43]~q ),
	.prn(vcc));
defparam \in_data_buffer[43] .is_wysiwyg = "true";
defparam \in_data_buffer[43] .power_up = "low";

dffeas \in_data_buffer[44] (
	.clk(wire_pll7_clk_0),
	.d(in_data[44]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[44]~q ),
	.prn(vcc));
defparam \in_data_buffer[44] .is_wysiwyg = "true";
defparam \in_data_buffer[44] .power_up = "low";

dffeas \in_data_buffer[45] (
	.clk(wire_pll7_clk_0),
	.d(in_data[45]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[45]~q ),
	.prn(vcc));
defparam \in_data_buffer[45] .is_wysiwyg = "true";
defparam \in_data_buffer[45] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~2_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut (
	clk,
	reset_n,
	dreg_0,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_0;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_1 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_avalon_st_handshake_clock_crosser_2 (
	wire_pll7_clk_0,
	W_alu_result_3,
	W_alu_result_2,
	r_sync_rst,
	uav_read,
	cp_valid,
	d_writedata_0,
	d_writedata_1,
	out_data_buffer_0,
	out_data_toggle_flopped,
	dreg_0,
	mem_used_1,
	out_data_buffer_65,
	out_data_buffer_38,
	out_data_buffer_39,
	altera_reset_synchronizer_int_chain_out,
	src_channel_12,
	Equal5,
	take_in_data,
	rst1,
	out_data_buffer_66,
	out_data_buffer_105,
	out_data_buffer_64,
	uav_write,
	Equal51,
	out_data_buffer_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	r_sync_rst;
input 	uav_read;
input 	cp_valid;
input 	d_writedata_0;
input 	d_writedata_1;
output 	out_data_buffer_0;
output 	out_data_toggle_flopped;
output 	dreg_0;
input 	mem_used_1;
output 	out_data_buffer_65;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_channel_12;
input 	Equal5;
output 	take_in_data;
input 	rst1;
output 	out_data_buffer_66;
output 	out_data_buffer_105;
output 	out_data_buffer_64;
input 	uav_write;
input 	Equal51;
output 	out_data_buffer_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_avalon_st_clock_crosser_1 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,uav_read,uav_write,uav_write,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,W_alu_result_3,W_alu_result_2,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_1,d_writedata_0}),
	.in_reset(r_sync_rst),
	.cp_valid(cp_valid),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.mem_used_1(mem_used_1),
	.out_data_buffer_65(out_data_buffer_65),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(out_data_buffer_39),
	.out_reset(altera_reset_synchronizer_int_chain_out),
	.src_channel_12(src_channel_12),
	.Equal5(Equal5),
	.take_in_data1(take_in_data),
	.rst1(rst1),
	.out_data_buffer_66(out_data_buffer_66),
	.out_data_buffer_105(out_data_buffer_105),
	.out_data_buffer_64(out_data_buffer_64),
	.Equal51(Equal51),
	.out_data_buffer_1(out_data_buffer_1),
	.clk_clk(clk_clk));

endmodule

module niosII_altera_avalon_st_clock_crosser_1 (
	wire_pll7_clk_0,
	in_data,
	in_reset,
	cp_valid,
	out_data_buffer_0,
	out_data_toggle_flopped1,
	dreg_0,
	mem_used_1,
	out_data_buffer_65,
	out_data_buffer_38,
	out_data_buffer_39,
	out_reset,
	src_channel_12,
	Equal5,
	take_in_data1,
	rst1,
	out_data_buffer_66,
	out_data_buffer_105,
	out_data_buffer_64,
	Equal51,
	out_data_buffer_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	[120:0] in_data;
input 	in_reset;
input 	cp_valid;
output 	out_data_buffer_0;
output 	out_data_toggle_flopped1;
output 	dreg_0;
input 	mem_used_1;
output 	out_data_buffer_65;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
input 	out_reset;
input 	src_channel_12;
input 	Equal5;
output 	take_in_data1;
input 	rst1;
output 	out_data_buffer_66;
output 	out_data_buffer_105;
output 	out_data_buffer_64;
input 	Equal51;
output 	out_data_buffer_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_to_in_synchronizer|dreg[0]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_toggle~q ;
wire \take_in_data~combout ;
wire \in_data_buffer[0]~q ;
wire \out_data_toggle_flopped~0_combout ;
wire \in_data_buffer[65]~q ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[39]~q ;
wire \in_data_buffer[66]~q ;
wire \in_data_buffer[105]~q ;
wire \in_data_buffer[64]~q ;
wire \in_data_buffer[1]~q ;


niosII_altera_std_synchronizer_nocut_3 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(\out_to_in_synchronizer|dreg[0]~q ));

niosII_altera_std_synchronizer_nocut_2 in_to_out_synchronizer(
	.dreg_0(dreg_0),
	.reset_n(out_reset),
	.din(\in_data_toggle~q ),
	.clk(clk_clk));

dffeas \out_data_buffer[0] (
	.clk(clk_clk),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas out_data_toggle_flopped(
	.clk(clk_clk),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

dffeas \out_data_buffer[65] (
	.clk(clk_clk),
	.d(\in_data_buffer[65]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_65),
	.prn(vcc));
defparam \out_data_buffer[65] .is_wysiwyg = "true";
defparam \out_data_buffer[65] .power_up = "low";

dffeas \out_data_buffer[38] (
	.clk(clk_clk),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[39] (
	.clk(clk_clk),
	.d(\in_data_buffer[39]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_39),
	.prn(vcc));
defparam \out_data_buffer[39] .is_wysiwyg = "true";
defparam \out_data_buffer[39] .power_up = "low";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(Equal5),
	.datab(src_channel_12),
	.datac(\in_data_toggle~q ),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(take_in_data1),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hEFFE;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \out_data_buffer[66] (
	.clk(clk_clk),
	.d(\in_data_buffer[66]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_66),
	.prn(vcc));
defparam \out_data_buffer[66] .is_wysiwyg = "true";
defparam \out_data_buffer[66] .power_up = "low";

dffeas \out_data_buffer[105] (
	.clk(clk_clk),
	.d(\in_data_buffer[105]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_105),
	.prn(vcc));
defparam \out_data_buffer[105] .is_wysiwyg = "true";
defparam \out_data_buffer[105] .power_up = "low";

dffeas \out_data_buffer[64] (
	.clk(clk_clk),
	.d(\in_data_buffer[64]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_64),
	.prn(vcc));
defparam \out_data_buffer[64] .is_wysiwyg = "true";
defparam \out_data_buffer[64] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(clk_clk),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(gnd),
	.datab(\in_data_toggle~q ),
	.datac(cp_valid),
	.datad(take_in_data1),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hC33C;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_data_toggle~q ),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb take_in_data(
	.dataa(cp_valid),
	.datab(Equal51),
	.datac(\in_data_toggle~q ),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hEFFE;
defparam take_in_data.sum_lutc_input = "datac";

dffeas \in_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(out_data_toggle_flopped1),
	.datab(dreg_0),
	.datac(rst1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[65] (
	.clk(wire_pll7_clk_0),
	.d(in_data[65]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[65]~q ),
	.prn(vcc));
defparam \in_data_buffer[65] .is_wysiwyg = "true";
defparam \in_data_buffer[65] .power_up = "low";

dffeas \in_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[39] (
	.clk(wire_pll7_clk_0),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[39]~q ),
	.prn(vcc));
defparam \in_data_buffer[39] .is_wysiwyg = "true";
defparam \in_data_buffer[39] .power_up = "low";

dffeas \in_data_buffer[66] (
	.clk(wire_pll7_clk_0),
	.d(in_data[66]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[66]~q ),
	.prn(vcc));
defparam \in_data_buffer[66] .is_wysiwyg = "true";
defparam \in_data_buffer[66] .power_up = "low";

dffeas \in_data_buffer[105] (
	.clk(wire_pll7_clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[105]~q ),
	.prn(vcc));
defparam \in_data_buffer[105] .is_wysiwyg = "true";
defparam \in_data_buffer[105] .power_up = "low";

dffeas \in_data_buffer[64] (
	.clk(wire_pll7_clk_0),
	.d(in_data[65]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[64]~q ),
	.prn(vcc));
defparam \in_data_buffer[64] .is_wysiwyg = "true";
defparam \in_data_buffer[64] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_2 (
	dreg_0,
	reset_n,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	reset_n;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_3 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_avalon_st_handshake_clock_crosser_3 (
	wire_pll7_clk_0,
	r_sync_rst,
	r_sync_rst1,
	saved_grant_1,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	hold_waitrequest,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	last_cycle,
	out_data_buffer_105,
	out_data_buffer_46,
	i_read,
	read_accepted,
	cp_valid,
	Equal1,
	uav_read,
	F_pc_8,
	F_pc_9,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	out_data_buffer_66,
	take_in_data,
	out_data_buffer_84,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	r_sync_rst1;
input 	saved_grant_1;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
input 	hold_waitrequest;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	out_valid;
input 	last_cycle;
output 	out_data_buffer_105;
output 	out_data_buffer_46;
input 	i_read;
input 	read_accepted;
input 	cp_valid;
input 	Equal1;
input 	uav_read;
input 	F_pc_8;
input 	F_pc_9;
input 	F_pc_0;
input 	F_pc_1;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_7;
output 	out_data_buffer_66;
output 	take_in_data;
output 	out_data_buffer_84;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_avalon_st_clock_crosser_2 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.in_reset(r_sync_rst),
	.out_reset(r_sync_rst1),
	.saved_grant_1(saved_grant_1),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(out_data_buffer_39),
	.out_data_buffer_40(out_data_buffer_40),
	.hold_waitrequest(hold_waitrequest),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid),
	.last_cycle(last_cycle),
	.out_data_buffer_105(out_data_buffer_105),
	.out_data_buffer_46(out_data_buffer_46),
	.i_read(i_read),
	.read_accepted(read_accepted),
	.cp_valid(cp_valid),
	.Equal1(Equal1),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,uav_read,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,F_pc_8,F_pc_7,F_pc_6,F_pc_5,
F_pc_4,F_pc_3,F_pc_2,F_pc_1,F_pc_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.F_pc_9(F_pc_9),
	.out_data_buffer_66(out_data_buffer_66),
	.take_in_data1(take_in_data),
	.out_data_buffer_84(out_data_buffer_84),
	.out_data_buffer_41(out_data_buffer_41),
	.out_data_buffer_42(out_data_buffer_42),
	.out_data_buffer_43(out_data_buffer_43),
	.out_data_buffer_44(out_data_buffer_44),
	.out_data_buffer_45(out_data_buffer_45));

endmodule

module niosII_altera_avalon_st_clock_crosser_2 (
	wire_pll7_clk_0,
	in_reset,
	out_reset,
	saved_grant_1,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	hold_waitrequest,
	out_data_toggle_flopped1,
	dreg_0,
	out_valid1,
	last_cycle,
	out_data_buffer_105,
	out_data_buffer_46,
	i_read,
	read_accepted,
	cp_valid,
	Equal1,
	in_data,
	F_pc_9,
	out_data_buffer_66,
	take_in_data1,
	out_data_buffer_84,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	in_reset;
input 	out_reset;
input 	saved_grant_1;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
input 	hold_waitrequest;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	out_valid1;
input 	last_cycle;
output 	out_data_buffer_105;
output 	out_data_buffer_46;
input 	i_read;
input 	read_accepted;
input 	cp_valid;
input 	Equal1;
input 	[120:0] in_data;
input 	F_pc_9;
output 	out_data_buffer_66;
output 	take_in_data1;
output 	out_data_buffer_84;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_to_in_synchronizer|dreg[0]~q ;
wire \take_in_data~combout ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[39]~q ;
wire \in_data_buffer[40]~q ;
wire \out_data_toggle_flopped~0_combout ;
wire \in_data_buffer[105]~q ;
wire \in_data_buffer[46]~q ;
wire \in_data_buffer[66]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_toggle~q ;
wire \in_data_buffer[84]~q ;
wire \in_data_buffer[41]~q ;
wire \in_data_buffer[42]~q ;
wire \in_data_buffer[43]~q ;
wire \in_data_buffer[44]~q ;
wire \in_data_buffer[45]~q ;


niosII_altera_std_synchronizer_nocut_5 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(\out_to_in_synchronizer|dreg[0]~q ));

niosII_altera_std_synchronizer_nocut_4 in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.dreg_0(dreg_0),
	.din(\in_data_toggle~q ));

dffeas \out_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[39] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[39]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_39),
	.prn(vcc));
defparam \out_data_buffer[39] .is_wysiwyg = "true";
defparam \out_data_buffer[39] .power_up = "low";

dffeas \out_data_buffer[40] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[40]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_40),
	.prn(vcc));
defparam \out_data_buffer[40] .is_wysiwyg = "true";
defparam \out_data_buffer[40] .power_up = "low";

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[105] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[105]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_105),
	.prn(vcc));
defparam \out_data_buffer[105] .is_wysiwyg = "true";
defparam \out_data_buffer[105] .power_up = "low";

dffeas \out_data_buffer[46] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[46]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_46),
	.prn(vcc));
defparam \out_data_buffer[46] .is_wysiwyg = "true";
defparam \out_data_buffer[46] .power_up = "low";

dffeas \out_data_buffer[66] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[66]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_66),
	.prn(vcc));
defparam \out_data_buffer[66] .is_wysiwyg = "true";
defparam \out_data_buffer[66] .power_up = "low";

cycloneive_lcell_comb \take_in_data~2 (
	.dataa(Equal1),
	.datab(\in_data_toggle~q ),
	.datac(\out_to_in_synchronizer|dreg[0]~q ),
	.datad(F_pc_9),
	.cin(gnd),
	.combout(take_in_data1),
	.cout());
defparam \take_in_data~2 .lut_mask = 16'hBEFF;
defparam \take_in_data~2 .sum_lutc_input = "datac";

dffeas \out_data_buffer[84] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[84]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_84),
	.prn(vcc));
defparam \out_data_buffer[84] .is_wysiwyg = "true";
defparam \out_data_buffer[84] .power_up = "low";

dffeas \out_data_buffer[41] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[41]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_41),
	.prn(vcc));
defparam \out_data_buffer[41] .is_wysiwyg = "true";
defparam \out_data_buffer[41] .power_up = "low";

dffeas \out_data_buffer[42] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[42]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_42),
	.prn(vcc));
defparam \out_data_buffer[42] .is_wysiwyg = "true";
defparam \out_data_buffer[42] .power_up = "low";

dffeas \out_data_buffer[43] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[43]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_43),
	.prn(vcc));
defparam \out_data_buffer[43] .is_wysiwyg = "true";
defparam \out_data_buffer[43] .power_up = "low";

dffeas \out_data_buffer[44] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[44]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_44),
	.prn(vcc));
defparam \out_data_buffer[44] .is_wysiwyg = "true";
defparam \out_data_buffer[44] .power_up = "low";

dffeas \out_data_buffer[45] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[45]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_45),
	.prn(vcc));
defparam \out_data_buffer[45] .is_wysiwyg = "true";
defparam \out_data_buffer[45] .power_up = "low";

cycloneive_lcell_comb take_in_data(
	.dataa(i_read),
	.datab(read_accepted),
	.datac(hold_waitrequest),
	.datad(take_in_data1),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hFFF7;
defparam take_in_data.sum_lutc_input = "datac";

dffeas \in_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[39] (
	.clk(wire_pll7_clk_0),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[39]~q ),
	.prn(vcc));
defparam \in_data_buffer[39] .is_wysiwyg = "true";
defparam \in_data_buffer[39] .power_up = "low";

dffeas \in_data_buffer[40] (
	.clk(wire_pll7_clk_0),
	.d(in_data[40]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[40]~q ),
	.prn(vcc));
defparam \in_data_buffer[40] .is_wysiwyg = "true";
defparam \in_data_buffer[40] .power_up = "low";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(dreg_0),
	.datab(out_data_toggle_flopped1),
	.datac(saved_grant_1),
	.datad(last_cycle),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[105] (
	.clk(wire_pll7_clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[105]~q ),
	.prn(vcc));
defparam \in_data_buffer[105] .is_wysiwyg = "true";
defparam \in_data_buffer[105] .power_up = "low";

dffeas \in_data_buffer[46] (
	.clk(wire_pll7_clk_0),
	.d(in_data[46]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[46]~q ),
	.prn(vcc));
defparam \in_data_buffer[46] .is_wysiwyg = "true";
defparam \in_data_buffer[46] .power_up = "low";

dffeas \in_data_buffer[66] (
	.clk(wire_pll7_clk_0),
	.d(in_data[66]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[66]~q ),
	.prn(vcc));
defparam \in_data_buffer[66] .is_wysiwyg = "true";
defparam \in_data_buffer[66] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(gnd),
	.datab(\in_data_toggle~q ),
	.datac(cp_valid),
	.datad(take_in_data1),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hC33C;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_data_toggle~q ),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

dffeas \in_data_buffer[84] (
	.clk(wire_pll7_clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[84]~q ),
	.prn(vcc));
defparam \in_data_buffer[84] .is_wysiwyg = "true";
defparam \in_data_buffer[84] .power_up = "low";

dffeas \in_data_buffer[41] (
	.clk(wire_pll7_clk_0),
	.d(in_data[41]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[41]~q ),
	.prn(vcc));
defparam \in_data_buffer[41] .is_wysiwyg = "true";
defparam \in_data_buffer[41] .power_up = "low";

dffeas \in_data_buffer[42] (
	.clk(wire_pll7_clk_0),
	.d(in_data[42]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[42]~q ),
	.prn(vcc));
defparam \in_data_buffer[42] .is_wysiwyg = "true";
defparam \in_data_buffer[42] .power_up = "low";

dffeas \in_data_buffer[43] (
	.clk(wire_pll7_clk_0),
	.d(in_data[43]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[43]~q ),
	.prn(vcc));
defparam \in_data_buffer[43] .is_wysiwyg = "true";
defparam \in_data_buffer[43] .power_up = "low";

dffeas \in_data_buffer[44] (
	.clk(wire_pll7_clk_0),
	.d(in_data[44]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[44]~q ),
	.prn(vcc));
defparam \in_data_buffer[44] .is_wysiwyg = "true";
defparam \in_data_buffer[44] .power_up = "low";

dffeas \in_data_buffer[45] (
	.clk(wire_pll7_clk_0),
	.d(in_data[45]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[45]~q ),
	.prn(vcc));
defparam \in_data_buffer[45] .is_wysiwyg = "true";
defparam \in_data_buffer[45] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_4 (
	clk,
	reset_n,
	dreg_0,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_0;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_5 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_avalon_st_handshake_clock_crosser_4 (
	wire_pll7_clk_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	out_data_toggle_flopped,
	dreg_0,
	in_data_toggle,
	out_valid,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	rp_valid,
	dreg_01,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_16,
	out_data_buffer_15,
	out_data_buffer_14,
	out_data_buffer_13,
	out_data_buffer_12,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	in_ready,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_22,
	out_data_21,
	out_data_20,
	out_data_19,
	out_data_18,
	out_data_17,
	out_data_16,
	out_data_15,
	out_data_14,
	out_data_13,
	out_data_12,
	out_data_10,
	out_data_9,
	out_data_8,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	in_data_toggle;
output 	out_valid;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
input 	rp_valid;
output 	dreg_01;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_16;
output 	out_data_buffer_15;
output 	out_data_buffer_14;
output 	out_data_buffer_13;
output 	out_data_buffer_12;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
output 	in_ready;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
input 	out_data_5;
input 	out_data_6;
input 	out_data_7;
input 	out_data_22;
input 	out_data_21;
input 	out_data_20;
input 	out_data_19;
input 	out_data_18;
input 	out_data_17;
input 	out_data_16;
input 	out_data_15;
input 	out_data_14;
input 	out_data_13;
input 	out_data_12;
input 	out_data_10;
input 	out_data_9;
input 	out_data_8;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_avalon_st_clock_crosser_3 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.out_reset(r_sync_rst),
	.in_reset(altera_reset_synchronizer_int_chain_out),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.in_data_toggle1(in_data_toggle),
	.out_valid1(out_valid),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_7(out_data_buffer_7),
	.rp_valid(rp_valid),
	.dreg_01(dreg_01),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_8(out_data_buffer_8),
	.in_ready(in_ready),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,out_data_22,out_data_21,out_data_20,out_data_19,out_data_18,out_data_17,out_data_16,out_data_15,out_data_14,out_data_13,out_data_12,gnd,out_data_10,out_data_9,out_data_8,out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,
out_data_1,out_data_0}),
	.clk_clk(clk_clk));

endmodule

module niosII_altera_avalon_st_clock_crosser_3 (
	wire_pll7_clk_0,
	out_reset,
	in_reset,
	out_data_toggle_flopped1,
	dreg_0,
	in_data_toggle1,
	out_valid1,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	rp_valid,
	dreg_01,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_16,
	out_data_buffer_15,
	out_data_buffer_14,
	out_data_buffer_13,
	out_data_buffer_12,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	in_ready,
	in_data,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	out_reset;
input 	in_reset;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	in_data_toggle1;
output 	out_valid1;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
input 	rp_valid;
output 	dreg_01;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_16;
output 	out_data_buffer_15;
output 	out_data_buffer_14;
output 	out_data_buffer_13;
output 	out_data_buffer_12;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
output 	in_ready;
input 	[120:0] in_data;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \in_data_toggle~0_combout ;
wire \take_in_data~combout ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[8]~q ;


niosII_altera_std_synchronizer_nocut_7 out_to_in_synchronizer(
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(dreg_01),
	.clk(clk_clk));

niosII_altera_std_synchronizer_nocut_6 in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.dreg_0(dreg_0),
	.din(in_data_toggle1));

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(dreg_0),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

dffeas in_data_toggle(
	.clk(clk_clk),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

cycloneive_lcell_comb \in_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(in_data_toggle1),
	.datad(dreg_01),
	.cin(gnd),
	.combout(in_ready),
	.cout());
defparam \in_ready~0 .lut_mask = 16'h0FF0;
defparam \in_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(gnd),
	.datac(rp_valid),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hA0AF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb take_in_data(
	.dataa(in_data_toggle1),
	.datab(dreg_01),
	.datac(rp_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hF6F6;
defparam take_in_data.sum_lutc_input = "datac";

dffeas \in_data_buffer[0] (
	.clk(clk_clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(clk_clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(clk_clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(clk_clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(clk_clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(clk_clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(clk_clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(clk_clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(clk_clk),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(clk_clk),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(clk_clk),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(clk_clk),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(clk_clk),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(clk_clk),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(clk_clk),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(clk_clk),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(clk_clk),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(clk_clk),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(clk_clk),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(clk_clk),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(clk_clk),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(clk_clk),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_6 (
	clk,
	reset_n,
	dreg_0,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_0;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_7 (
	reset_n,
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_avalon_st_handshake_clock_crosser_5 (
	wire_pll7_clk_0,
	r_sync_rst,
	r_sync_rst1,
	out_data_toggle_flopped,
	dreg_0,
	in_data_toggle,
	dreg_01,
	take_in_data,
	rp_valid,
	out_valid,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_16,
	out_data_buffer_15,
	out_data_buffer_14,
	out_data_buffer_13,
	out_data_buffer_12,
	out_data_buffer_11,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_buffer_27,
	out_data_buffer_28,
	out_data_buffer_29,
	out_data_buffer_30,
	out_data_buffer_31,
	out_data_11,
	out_data_13,
	out_data_16,
	out_data_12,
	out_data_5,
	out_data_14,
	out_data_15,
	out_data_10,
	out_data_9,
	out_data_8,
	out_data_7,
	out_data_6,
	out_data_21,
	out_data_30,
	out_data_29,
	out_data_28,
	out_data_27,
	out_data_26,
	out_data_25,
	out_data_24,
	out_data_23,
	out_data_22,
	out_data_20,
	out_data_19,
	out_data_18,
	out_data_17,
	out_data_31)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	r_sync_rst1;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	in_data_toggle;
output 	dreg_01;
input 	take_in_data;
input 	rp_valid;
output 	out_valid;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_16;
output 	out_data_buffer_15;
output 	out_data_buffer_14;
output 	out_data_buffer_13;
output 	out_data_buffer_12;
output 	out_data_buffer_11;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
output 	out_data_buffer_27;
output 	out_data_buffer_28;
output 	out_data_buffer_29;
output 	out_data_buffer_30;
output 	out_data_buffer_31;
input 	out_data_11;
input 	out_data_13;
input 	out_data_16;
input 	out_data_12;
input 	out_data_5;
input 	out_data_14;
input 	out_data_15;
input 	out_data_10;
input 	out_data_9;
input 	out_data_8;
input 	out_data_7;
input 	out_data_6;
input 	out_data_21;
input 	out_data_30;
input 	out_data_29;
input 	out_data_28;
input 	out_data_27;
input 	out_data_26;
input 	out_data_25;
input 	out_data_24;
input 	out_data_23;
input 	out_data_22;
input 	out_data_20;
input 	out_data_19;
input 	out_data_18;
input 	out_data_17;
input 	out_data_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_avalon_st_clock_crosser_4 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.out_reset(r_sync_rst),
	.in_reset(r_sync_rst1),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.in_data_toggle1(in_data_toggle),
	.dreg_01(dreg_01),
	.take_in_data(take_in_data),
	.rp_valid(rp_valid),
	.out_valid1(out_valid),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_8(out_data_buffer_8),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,out_data_31,out_data_30,out_data_29,out_data_28,out_data_27,out_data_26,out_data_25,out_data_24,out_data_23,out_data_22,out_data_21,out_data_20,out_data_19,out_data_18,out_data_17,out_data_16,out_data_15,out_data_14,out_data_13,out_data_12,out_data_11,out_data_10,
out_data_9,out_data_8,out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,out_data_1,out_data_0}),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_31(out_data_buffer_31));

endmodule

module niosII_altera_avalon_st_clock_crosser_4 (
	wire_pll7_clk_0,
	out_reset,
	in_reset,
	out_data_toggle_flopped1,
	dreg_0,
	in_data_toggle1,
	dreg_01,
	take_in_data,
	rp_valid,
	out_valid1,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_16,
	out_data_buffer_15,
	out_data_buffer_14,
	out_data_buffer_13,
	out_data_buffer_12,
	out_data_buffer_11,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	in_data,
	out_data_buffer_27,
	out_data_buffer_28,
	out_data_buffer_29,
	out_data_buffer_30,
	out_data_buffer_31)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	out_reset;
input 	in_reset;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	in_data_toggle1;
output 	dreg_01;
input 	take_in_data;
input 	rp_valid;
output 	out_valid1;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_16;
output 	out_data_buffer_15;
output 	out_data_buffer_14;
output 	out_data_buffer_13;
output 	out_data_buffer_12;
output 	out_data_buffer_11;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
input 	[120:0] in_data;
output 	out_data_buffer_27;
output 	out_data_buffer_28;
output 	out_data_buffer_29;
output 	out_data_buffer_30;
output 	out_data_buffer_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \in_data_toggle~0_combout ;
wire \take_in_data~0_combout ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[29]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[31]~q ;


niosII_altera_std_synchronizer_nocut_9 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(dreg_01));

niosII_altera_std_synchronizer_nocut_8 in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.dreg_0(dreg_0),
	.din(in_data_toggle1));

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(dreg_0),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(take_in_data),
	.datac(rp_valid),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(rp_valid),
	.datab(in_data_toggle1),
	.datac(dreg_01),
	.datad(take_in_data),
	.cin(gnd),
	.combout(\take_in_data~0_combout ),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hBEFF;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_8 (
	clk,
	reset_n,
	dreg_0,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_0;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_9 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_avalon_st_handshake_clock_crosser_6 (
	wire_pll7_clk_0,
	r_sync_rst,
	r_sync_rst1,
	mem_84_0,
	mem_66_0,
	in_data_toggle,
	dreg_0,
	take_in_data,
	out_data_toggle_flopped,
	dreg_01,
	rp_valid,
	out_valid,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_16,
	out_data_buffer_12,
	out_data_buffer_5,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_21,
	out_data_buffer_30,
	out_data_buffer_29,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_31,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_11,
	out_data_13,
	out_data_16,
	out_data_12,
	out_data_5,
	out_data_14,
	out_data_15,
	out_data_10,
	out_data_9,
	out_data_8,
	out_data_7,
	out_data_6,
	out_data_21,
	out_data_30,
	out_data_29,
	out_data_28,
	out_data_27,
	out_data_26,
	out_data_25,
	out_data_24,
	out_data_23,
	out_data_22,
	out_data_20,
	out_data_19,
	out_data_18,
	out_data_17,
	out_data_31)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	r_sync_rst1;
input 	mem_84_0;
input 	mem_66_0;
output 	in_data_toggle;
output 	dreg_0;
output 	take_in_data;
output 	out_data_toggle_flopped;
output 	dreg_01;
input 	rp_valid;
output 	out_valid;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_16;
output 	out_data_buffer_12;
output 	out_data_buffer_5;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_21;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_31;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
input 	out_data_11;
input 	out_data_13;
input 	out_data_16;
input 	out_data_12;
input 	out_data_5;
input 	out_data_14;
input 	out_data_15;
input 	out_data_10;
input 	out_data_9;
input 	out_data_8;
input 	out_data_7;
input 	out_data_6;
input 	out_data_21;
input 	out_data_30;
input 	out_data_29;
input 	out_data_28;
input 	out_data_27;
input 	out_data_26;
input 	out_data_25;
input 	out_data_24;
input 	out_data_23;
input 	out_data_22;
input 	out_data_20;
input 	out_data_19;
input 	out_data_18;
input 	out_data_17;
input 	out_data_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_avalon_st_clock_crosser_5 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.out_reset(r_sync_rst),
	.in_reset(r_sync_rst1),
	.mem_84_0(mem_84_0),
	.mem_66_0(mem_66_0),
	.in_data_toggle1(in_data_toggle),
	.dreg_0(dreg_0),
	.take_in_data(take_in_data),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_01(dreg_01),
	.rp_valid(rp_valid),
	.out_valid1(out_valid),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_31(out_data_buffer_31),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,out_data_31,out_data_30,out_data_29,out_data_28,out_data_27,out_data_26,out_data_25,out_data_24,out_data_23,out_data_22,out_data_21,out_data_20,out_data_19,out_data_18,out_data_17,out_data_16,out_data_15,out_data_14,out_data_13,out_data_12,out_data_11,out_data_10,
out_data_9,out_data_8,out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,out_data_1,out_data_0}));

endmodule

module niosII_altera_avalon_st_clock_crosser_5 (
	wire_pll7_clk_0,
	out_reset,
	in_reset,
	mem_84_0,
	mem_66_0,
	in_data_toggle1,
	dreg_0,
	take_in_data,
	out_data_toggle_flopped1,
	dreg_01,
	rp_valid,
	out_valid1,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_16,
	out_data_buffer_12,
	out_data_buffer_5,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_21,
	out_data_buffer_30,
	out_data_buffer_29,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_31,
	in_data)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	out_reset;
input 	in_reset;
input 	mem_84_0;
input 	mem_66_0;
output 	in_data_toggle1;
output 	dreg_0;
output 	take_in_data;
output 	out_data_toggle_flopped1;
output 	dreg_01;
input 	rp_valid;
output 	out_valid1;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_16;
output 	out_data_buffer_12;
output 	out_data_buffer_5;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_21;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_31;
input 	[120:0] in_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \in_data_toggle~0_combout ;
wire \take_in_data~1_combout ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[29]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[31]~q ;


niosII_altera_std_synchronizer_nocut_11 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.dreg_0(dreg_0),
	.din(out_data_toggle_flopped1));

niosII_altera_std_synchronizer_nocut_10 in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.din(in_data_toggle1),
	.dreg_0(dreg_01));

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(mem_84_0),
	.datab(mem_66_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(take_in_data),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hEEEE;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(dreg_01),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_01),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(take_in_data),
	.datac(rp_valid),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_in_data~1 (
	.dataa(take_in_data),
	.datab(rp_valid),
	.datac(in_data_toggle1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\take_in_data~1_combout ),
	.cout());
defparam \take_in_data~1 .lut_mask = 16'hEFFE;
defparam \take_in_data~1 .sum_lutc_input = "datac";

dffeas \in_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_10 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_11 (
	clk,
	reset_n,
	dreg_0,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_0;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_avalon_st_handshake_clock_crosser_7 (
	wire_pll7_clk_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	out_data_toggle_flopped,
	dreg_0,
	in_ready,
	rp_valid,
	out_valid,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_0,
	out_data_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	in_ready;
input 	rp_valid;
output 	out_valid;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
input 	out_data_0;
input 	out_data_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_avalon_st_clock_crosser_6 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.out_reset(r_sync_rst),
	.in_reset(altera_reset_synchronizer_int_chain_out),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.in_ready(in_ready),
	.rp_valid(rp_valid),
	.out_valid1(out_valid),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,out_data_1,out_data_0}),
	.clk_clk(clk_clk));

endmodule

module niosII_altera_avalon_st_clock_crosser_6 (
	wire_pll7_clk_0,
	out_reset,
	in_reset,
	out_data_toggle_flopped1,
	dreg_0,
	in_ready,
	rp_valid,
	out_valid1,
	out_data_buffer_0,
	out_data_buffer_1,
	in_data,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	out_reset;
input 	in_reset;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	in_ready;
input 	rp_valid;
output 	out_valid1;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
input 	[120:0] in_data;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_to_in_synchronizer|dreg[0]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_toggle~q ;
wire \take_in_data~combout ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;


niosII_altera_std_synchronizer_nocut_13 out_to_in_synchronizer(
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(\out_to_in_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

niosII_altera_std_synchronizer_nocut_12 in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.dreg_0(dreg_0),
	.din(\in_data_toggle~q ));

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(dreg_0),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb \in_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_data_toggle~q ),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(in_ready),
	.cout());
defparam \in_ready~0 .lut_mask = 16'h0FF0;
defparam \in_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(\in_data_toggle~q ),
	.datab(gnd),
	.datac(rp_valid),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hA0AF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(clk_clk),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_data_toggle~q ),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb take_in_data(
	.dataa(\in_data_toggle~q ),
	.datab(\out_to_in_synchronizer|dreg[0]~q ),
	.datac(rp_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hF6F6;
defparam take_in_data.sum_lutc_input = "datac";

dffeas \in_data_buffer[0] (
	.clk(clk_clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(clk_clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_12 (
	clk,
	reset_n,
	dreg_0,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_0;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_13 (
	reset_n,
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_avalon_st_clock_crosser_7 (
	wire_pll7_clk_0,
	in_data,
	in_reset,
	cp_valid,
	out_reset,
	Equal13,
	in_data_toggle1,
	dreg_0,
	out_data_toggle_flopped1,
	dreg_01,
	av_waitrequest,
	mem_used_1,
	out_data_buffer_66,
	out_data_buffer_38,
	out_data_buffer_7,
	out_data_buffer_65,
	out_data_buffer_105,
	out_data_buffer_64,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_10,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	[120:0] in_data;
input 	in_reset;
input 	cp_valid;
input 	out_reset;
input 	Equal13;
output 	in_data_toggle1;
output 	dreg_0;
output 	out_data_toggle_flopped1;
output 	dreg_01;
input 	av_waitrequest;
input 	mem_used_1;
output 	out_data_buffer_66;
output 	out_data_buffer_38;
output 	out_data_buffer_7;
output 	out_data_buffer_65;
output 	out_data_buffer_105;
output 	out_data_buffer_64;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_10;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \in_data_toggle~0_combout ;
wire \out_data_toggle_flopped~0_combout ;
wire \take_in_data~combout ;
wire \in_data_buffer[66]~q ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[65]~q ;
wire \in_data_buffer[105]~q ;
wire \in_data_buffer[64]~q ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[6]~q ;


niosII_altera_std_synchronizer_nocut_15 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.dreg_0(dreg_0),
	.din(out_data_toggle_flopped1));

niosII_altera_std_synchronizer_nocut_14 in_to_out_synchronizer(
	.reset_n(out_reset),
	.din(in_data_toggle1),
	.dreg_0(dreg_01),
	.clk(clk_clk));

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

dffeas out_data_toggle_flopped(
	.clk(clk_clk),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

dffeas \out_data_buffer[66] (
	.clk(clk_clk),
	.d(\in_data_buffer[66]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_66),
	.prn(vcc));
defparam \out_data_buffer[66] .is_wysiwyg = "true";
defparam \out_data_buffer[66] .power_up = "low";

dffeas \out_data_buffer[38] (
	.clk(clk_clk),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(clk_clk),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[65] (
	.clk(clk_clk),
	.d(\in_data_buffer[65]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_65),
	.prn(vcc));
defparam \out_data_buffer[65] .is_wysiwyg = "true";
defparam \out_data_buffer[65] .power_up = "low";

dffeas \out_data_buffer[105] (
	.clk(clk_clk),
	.d(\in_data_buffer[105]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_105),
	.prn(vcc));
defparam \out_data_buffer[105] .is_wysiwyg = "true";
defparam \out_data_buffer[105] .power_up = "low";

dffeas \out_data_buffer[64] (
	.clk(clk_clk),
	.d(\in_data_buffer[64]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_64),
	.prn(vcc));
defparam \out_data_buffer[64] .is_wysiwyg = "true";
defparam \out_data_buffer[64] .power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(clk_clk),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(clk_clk),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(clk_clk),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(clk_clk),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(clk_clk),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(clk_clk),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(clk_clk),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(clk_clk),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(cp_valid),
	.datac(Equal13),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(out_data_toggle_flopped1),
	.datab(dreg_01),
	.datac(av_waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb take_in_data(
	.dataa(cp_valid),
	.datab(Equal13),
	.datac(in_data_toggle1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hEFFE;
defparam take_in_data.sum_lutc_input = "datac";

dffeas \in_data_buffer[66] (
	.clk(wire_pll7_clk_0),
	.d(in_data[66]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[66]~q ),
	.prn(vcc));
defparam \in_data_buffer[66] .is_wysiwyg = "true";
defparam \in_data_buffer[66] .power_up = "low";

dffeas \in_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[65] (
	.clk(wire_pll7_clk_0),
	.d(in_data[65]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[65]~q ),
	.prn(vcc));
defparam \in_data_buffer[65] .is_wysiwyg = "true";
defparam \in_data_buffer[65] .power_up = "low";

dffeas \in_data_buffer[105] (
	.clk(wire_pll7_clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[105]~q ),
	.prn(vcc));
defparam \in_data_buffer[105] .is_wysiwyg = "true";
defparam \in_data_buffer[105] .power_up = "low";

dffeas \in_data_buffer[64] (
	.clk(wire_pll7_clk_0),
	.d(in_data[65]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[64]~q ),
	.prn(vcc));
defparam \in_data_buffer[64] .is_wysiwyg = "true";
defparam \in_data_buffer[64] .power_up = "low";

dffeas \in_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_14 (
	reset_n,
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_std_synchronizer_nocut_15 (
	clk,
	reset_n,
	dreg_0,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_0;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosII_altera_merlin_master_agent (
	clk,
	r_sync_rst,
	uav_read,
	hold_waitrequest1,
	d_write,
	write_accepted,
	cp_valid)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	r_sync_rst;
input 	uav_read;
output 	hold_waitrequest1;
input 	d_write;
input 	write_accepted;
output 	cp_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas hold_waitrequest(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(hold_waitrequest1),
	.prn(vcc));
defparam hold_waitrequest.is_wysiwyg = "true";
defparam hold_waitrequest.power_up = "low";

cycloneive_lcell_comb \cp_valid~0 (
	.dataa(hold_waitrequest1),
	.datab(uav_read),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(cp_valid),
	.cout());
defparam \cp_valid~0 .lut_mask = 16'hFEFF;
defparam \cp_valid~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_master_agent_1 (
	hold_waitrequest,
	i_read,
	read_accepted,
	cp_valid1)/* synthesis synthesis_greybox=1 */;
input 	hold_waitrequest;
input 	i_read;
input 	read_accepted;
output 	cp_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb cp_valid(
	.dataa(hold_waitrequest),
	.datab(gnd),
	.datac(i_read),
	.datad(read_accepted),
	.cin(gnd),
	.combout(cp_valid1),
	.cout());
defparam cp_valid.lut_mask = 16'hAFFF;
defparam cp_valid.sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_master_translator (
	clk,
	reset,
	d_read,
	read_accepted1,
	uav_read,
	hold_waitrequest,
	d_write,
	write_accepted1,
	WideOr1,
	WideOr0,
	WideOr01,
	av_waitrequest,
	uav_write)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	d_read;
output 	read_accepted1;
output 	uav_read;
input 	hold_waitrequest;
input 	d_write;
output 	write_accepted1;
input 	WideOr1;
input 	WideOr0;
input 	WideOr01;
output 	av_waitrequest;
output 	uav_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;
wire \read_accepted~1_combout ;
wire \write_accepted~0_combout ;
wire \end_begintransfer~0_combout ;
wire \end_begintransfer~q ;
wire \av_waitrequest~0_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cycloneive_lcell_comb \uav_read~0 (
	.dataa(d_read),
	.datab(gnd),
	.datac(gnd),
	.datad(read_accepted1),
	.cin(gnd),
	.combout(uav_read),
	.cout());
defparam \uav_read~0 .lut_mask = 16'hAAFF;
defparam \uav_read~0 .sum_lutc_input = "datac";

dffeas write_accepted(
	.clk(clk),
	.d(\write_accepted~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(write_accepted1),
	.prn(vcc));
defparam write_accepted.is_wysiwyg = "true";
defparam write_accepted.power_up = "low";

cycloneive_lcell_comb \av_waitrequest~1 (
	.dataa(d_read),
	.datab(WideOr1),
	.datac(d_write),
	.datad(\av_waitrequest~0_combout ),
	.cin(gnd),
	.combout(av_waitrequest),
	.cout());
defparam \av_waitrequest~1 .lut_mask = 16'h8DFF;
defparam \av_waitrequest~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \uav_write~0 (
	.dataa(d_write),
	.datab(gnd),
	.datac(gnd),
	.datad(write_accepted1),
	.cin(gnd),
	.combout(uav_write),
	.cout());
defparam \uav_write~0 .lut_mask = 16'hAAFF;
defparam \uav_write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~0 (
	.dataa(hold_waitrequest),
	.datab(WideOr0),
	.datac(WideOr01),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_accepted~0_combout ),
	.cout());
defparam \read_accepted~0 .lut_mask = 16'hFEFE;
defparam \read_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~1 (
	.dataa(WideOr1),
	.datab(read_accepted1),
	.datac(d_read),
	.datad(\read_accepted~0_combout ),
	.cin(gnd),
	.combout(\read_accepted~1_combout ),
	.cout());
defparam \read_accepted~1 .lut_mask = 16'hFFFE;
defparam \read_accepted~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_accepted~0 (
	.dataa(av_waitrequest),
	.datab(write_accepted1),
	.datac(d_write),
	.datad(\read_accepted~0_combout ),
	.cin(gnd),
	.combout(\write_accepted~0_combout ),
	.cout());
defparam \write_accepted~0 .lut_mask = 16'hFFFE;
defparam \write_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \end_begintransfer~0 (
	.dataa(uav_write),
	.datab(uav_read),
	.datac(\end_begintransfer~q ),
	.datad(\read_accepted~0_combout ),
	.cin(gnd),
	.combout(\end_begintransfer~0_combout ),
	.cout());
defparam \end_begintransfer~0 .lut_mask = 16'hFEFF;
defparam \end_begintransfer~0 .sum_lutc_input = "datac";

dffeas end_begintransfer(
	.clk(clk),
	.d(\end_begintransfer~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\end_begintransfer~q ),
	.prn(vcc));
defparam end_begintransfer.is_wysiwyg = "true";
defparam end_begintransfer.power_up = "low";

cycloneive_lcell_comb \av_waitrequest~0 (
	.dataa(\end_begintransfer~q ),
	.datab(write_accepted1),
	.datac(\read_accepted~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_waitrequest~0_combout ),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hFEFE;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_master_translator_1 (
	clk,
	reset,
	hold_waitrequest,
	saved_grant_1,
	i_read,
	read_accepted1,
	Equal1,
	uav_read1,
	F_pc_9,
	last_cycle,
	waitrequest,
	mem_used_1,
	take_in_data,
	out_data_toggle_flopped,
	dreg_0,
	src1_valid,
	read_accepted2,
	src1_valid1,
	saved_grant_11)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	hold_waitrequest;
input 	saved_grant_1;
input 	i_read;
output 	read_accepted1;
input 	Equal1;
output 	uav_read1;
input 	F_pc_9;
input 	last_cycle;
input 	waitrequest;
input 	mem_used_1;
input 	take_in_data;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	src1_valid;
output 	read_accepted2;
input 	src1_valid1;
input 	saved_grant_11;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~6_combout ;
wire \read_accepted~3_combout ;
wire \read_accepted~4_combout ;
wire \read_accepted~5_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cycloneive_lcell_comb uav_read(
	.dataa(gnd),
	.datab(gnd),
	.datac(i_read),
	.datad(read_accepted1),
	.cin(gnd),
	.combout(uav_read1),
	.cout());
defparam uav_read.lut_mask = 16'h0FFF;
defparam uav_read.sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~2 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(gnd),
	.datad(src1_valid),
	.cin(gnd),
	.combout(read_accepted2),
	.cout());
defparam \read_accepted~2 .lut_mask = 16'h66FF;
defparam \read_accepted~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~6 (
	.dataa(waitrequest),
	.datab(mem_used_1),
	.datac(F_pc_9),
	.datad(saved_grant_11),
	.cin(gnd),
	.combout(\read_accepted~6_combout ),
	.cout());
defparam \read_accepted~6 .lut_mask = 16'hFFF7;
defparam \read_accepted~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~3 (
	.dataa(saved_grant_1),
	.datab(last_cycle),
	.datac(Equal1),
	.datad(\read_accepted~6_combout ),
	.cin(gnd),
	.combout(\read_accepted~3_combout ),
	.cout());
defparam \read_accepted~3 .lut_mask = 16'hFFAC;
defparam \read_accepted~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~4 (
	.dataa(hold_waitrequest),
	.datab(i_read),
	.datac(take_in_data),
	.datad(\read_accepted~3_combout ),
	.cin(gnd),
	.combout(\read_accepted~4_combout ),
	.cout());
defparam \read_accepted~4 .lut_mask = 16'hFFFB;
defparam \read_accepted~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~5 (
	.dataa(read_accepted2),
	.datab(read_accepted1),
	.datac(\read_accepted~4_combout ),
	.datad(src1_valid1),
	.cin(gnd),
	.combout(\read_accepted~5_combout ),
	.cout());
defparam \read_accepted~5 .lut_mask = 16'hFEFF;
defparam \read_accepted~5 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_agent (
	mem_used_1,
	uav_read,
	cp_valid,
	Equal3,
	m0_read1,
	m0_read2)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	uav_read;
input 	cp_valid;
input 	Equal3;
output 	m0_read1;
output 	m0_read2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb m0_read(
	.dataa(mem_used_1),
	.datab(uav_read),
	.datac(cp_valid),
	.datad(Equal3),
	.cin(gnd),
	.combout(m0_read1),
	.cout());
defparam m0_read.lut_mask = 16'hBFFF;
defparam m0_read.sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_read~0 (
	.dataa(Equal3),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(m0_read2),
	.cout());
defparam \m0_read~0 .lut_mask = 16'hAAFF;
defparam \m0_read~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_agent_1 (
	mem,
	WideOr1,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	mem;
input 	WideOr1;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \rf_source_valid~0 (
	.dataa(WideOr1),
	.datab(mem),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(rf_source_valid),
	.cout());
defparam \rf_source_valid~0 .lut_mask = 16'hEEEE;
defparam \rf_source_valid~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_agent_2 (
	src_payload_0,
	p1_wr_strobe,
	mem_used_0,
	mem_105_0,
	read_latency_shift_reg_0,
	mem_used_01,
	rp_valid1,
	WideOr0,
	rf_sink_ready,
	out_data_buffer_64,
	nonposted_write_endofpacket,
	rp_valid2,
	WideOr1)/* synthesis synthesis_greybox=1 */;
input 	src_payload_0;
input 	p1_wr_strobe;
input 	mem_used_0;
input 	mem_105_0;
input 	read_latency_shift_reg_0;
input 	mem_used_01;
output 	rp_valid1;
input 	WideOr0;
output 	rf_sink_ready;
input 	out_data_buffer_64;
output 	nonposted_write_endofpacket;
output 	rp_valid2;
input 	WideOr1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_merlin_burst_uncompressor_2 uncompressor(
	.mem_used_0(mem_used_0),
	.mem_105_0(mem_105_0),
	.rp_valid(rp_valid1),
	.WideOr0(WideOr0),
	.sink_ready(rf_sink_ready));

cycloneive_lcell_comb \rp_valid~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(rp_valid1),
	.cout());
defparam \rp_valid~0 .lut_mask = 16'h0FFF;
defparam \rp_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nonposted_write_endofpacket~0 (
	.dataa(WideOr1),
	.datab(src_payload_0),
	.datac(p1_wr_strobe),
	.datad(out_data_buffer_64),
	.cin(gnd),
	.combout(nonposted_write_endofpacket),
	.cout());
defparam \nonposted_write_endofpacket~0 .lut_mask = 16'hFEFF;
defparam \nonposted_write_endofpacket~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb rp_valid(
	.dataa(read_latency_shift_reg_0),
	.datab(mem_used_01),
	.datac(mem_used_0),
	.datad(mem_105_0),
	.cin(gnd),
	.combout(rp_valid2),
	.cout());
defparam rp_valid.lut_mask = 16'hFFFE;
defparam rp_valid.sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_burst_uncompressor_2 (
	mem_used_0,
	mem_105_0,
	rp_valid,
	WideOr0,
	sink_ready)/* synthesis synthesis_greybox=1 */;
input 	mem_used_0;
input 	mem_105_0;
input 	rp_valid;
input 	WideOr0;
output 	sink_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \sink_ready~0 (
	.dataa(mem_used_0),
	.datab(mem_105_0),
	.datac(rp_valid),
	.datad(WideOr0),
	.cin(gnd),
	.combout(sink_ready),
	.cout());
defparam \sink_ready~0 .lut_mask = 16'hEFFF;
defparam \sink_ready~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_agent_3 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_105_0,
	mem_used_01,
	rp_valid1,
	rp_valid2)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_105_0;
input 	mem_used_01;
output 	rp_valid1;
output 	rp_valid2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb rp_valid(
	.dataa(read_latency_shift_reg_0),
	.datab(mem_used_0),
	.datac(mem_105_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(rp_valid1),
	.cout());
defparam rp_valid.lut_mask = 16'hFFFE;
defparam rp_valid.sum_lutc_input = "datac";

cycloneive_lcell_comb \rp_valid~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(rp_valid2),
	.cout());
defparam \rp_valid~0 .lut_mask = 16'h0FFF;
defparam \rp_valid~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_agent_10 (
	wire_pll7_clk_0,
	byteen_reg_0,
	byteen_reg_1,
	r_sync_rst,
	entries_1,
	entries_0,
	d_write,
	write_accepted,
	d_byteenable_0,
	saved_grant_0,
	d_byteenable_1,
	use_reg,
	saved_grant_1,
	WideOr0,
	Equal0,
	Equal1,
	WideOr1,
	m0_write1,
	mem_used_7,
	src_data_66,
	src_valid,
	src12_valid,
	m0_write2,
	out_valid,
	mem_used_0,
	mem_87_0,
	rp_valid1,
	mem_54_0,
	burst_uncompress_address_base_1,
	burst_uncompress_address_offset_1,
	mem_19_0,
	comb,
	cp_ready1,
	mem_57_0,
	source_addr_1,
	cp_ready2,
	rf_source_data_87)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	byteen_reg_0;
input 	byteen_reg_1;
input 	r_sync_rst;
input 	entries_1;
input 	entries_0;
input 	d_write;
input 	write_accepted;
input 	d_byteenable_0;
input 	saved_grant_0;
input 	d_byteenable_1;
input 	use_reg;
input 	saved_grant_1;
output 	WideOr0;
input 	Equal0;
input 	Equal1;
input 	WideOr1;
output 	m0_write1;
input 	mem_used_7;
input 	src_data_66;
input 	src_valid;
input 	src12_valid;
output 	m0_write2;
input 	out_valid;
input 	mem_used_0;
input 	mem_87_0;
output 	rp_valid1;
input 	mem_54_0;
output 	burst_uncompress_address_base_1;
output 	burst_uncompress_address_offset_1;
input 	mem_19_0;
output 	comb;
output 	cp_ready1;
input 	mem_57_0;
output 	source_addr_1;
output 	cp_ready2;
output 	rf_source_data_87;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~0_combout ;
wire \WideOr0~1_combout ;
wire \m0_write~3_combout ;
wire \m0_write~4_combout ;


niosII_altera_merlin_burst_uncompressor_10 uncompressor(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.out_valid(out_valid),
	.mem_used_0(mem_used_0),
	.mem_87_0(mem_87_0),
	.mem_54_0(mem_54_0),
	.burst_uncompress_address_base_1(burst_uncompress_address_base_1),
	.burst_uncompress_address_offset_1(burst_uncompress_address_offset_1),
	.mem_19_0(mem_19_0),
	.comb(comb),
	.mem_57_0(mem_57_0),
	.source_addr_1(source_addr_1));

cycloneive_lcell_comb \WideOr0~2 (
	.dataa(\WideOr0~0_combout ),
	.datab(\WideOr0~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~2 .lut_mask = 16'hEEEE;
defparam \WideOr0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_write~2 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(m0_write1),
	.cout());
defparam \m0_write~2 .lut_mask = 16'hEEFF;
defparam \m0_write~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb m0_write(
	.dataa(src_valid),
	.datab(src12_valid),
	.datac(Equal1),
	.datad(\m0_write~4_combout ),
	.cin(gnd),
	.combout(m0_write2),
	.cout());
defparam m0_write.lut_mask = 16'hF7FF;
defparam m0_write.sum_lutc_input = "datac";

cycloneive_lcell_comb rp_valid(
	.dataa(out_valid),
	.datab(mem_used_0),
	.datac(mem_87_0),
	.datad(gnd),
	.cin(gnd),
	.combout(rp_valid1),
	.cout());
defparam rp_valid.lut_mask = 16'hFEFE;
defparam rp_valid.sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~0 (
	.dataa(gnd),
	.datab(mem_87_0),
	.datac(out_valid),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(comb),
	.cout());
defparam \comb~0 .lut_mask = 16'hFFFC;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb cp_ready(
	.dataa(mem_used_7),
	.datab(Equal0),
	.datac(\WideOr0~0_combout ),
	.datad(\WideOr0~1_combout ),
	.cin(gnd),
	.combout(cp_ready1),
	.cout());
defparam cp_ready.lut_mask = 16'hFFFE;
defparam cp_ready.sum_lutc_input = "datac";

cycloneive_lcell_comb \cp_ready~2 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\WideOr0~0_combout ),
	.datad(\WideOr0~1_combout ),
	.cin(gnd),
	.combout(cp_ready2),
	.cout());
defparam \cp_ready~2 .lut_mask = 16'hFFFB;
defparam \cp_ready~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rf_source_data[87]~2 (
	.dataa(\WideOr0~0_combout ),
	.datab(\WideOr0~1_combout ),
	.datac(src_data_66),
	.datad(WideOr1),
	.cin(gnd),
	.combout(rf_source_data_87),
	.cout());
defparam \rf_source_data[87]~2 .lut_mask = 16'hFFF7;
defparam \rf_source_data[87]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(saved_grant_0),
	.datab(d_byteenable_0),
	.datac(d_byteenable_1),
	.datad(use_reg),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hFEFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~1 (
	.dataa(saved_grant_1),
	.datab(use_reg),
	.datac(byteen_reg_0),
	.datad(byteen_reg_1),
	.cin(gnd),
	.combout(\WideOr0~1_combout ),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hFFB8;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_write~3 (
	.dataa(mem_used_7),
	.datab(saved_grant_0),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\m0_write~3_combout ),
	.cout());
defparam \m0_write~3 .lut_mask = 16'hFDFF;
defparam \m0_write~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_write~4 (
	.dataa(\WideOr0~0_combout ),
	.datab(\WideOr0~1_combout ),
	.datac(\m0_write~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\m0_write~4_combout ),
	.cout());
defparam \m0_write~4 .lut_mask = 16'hFEFE;
defparam \m0_write~4 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_burst_uncompressor_10 (
	clk,
	reset,
	out_valid,
	mem_used_0,
	mem_87_0,
	mem_54_0,
	burst_uncompress_address_base_1,
	burst_uncompress_address_offset_1,
	mem_19_0,
	comb,
	mem_57_0,
	source_addr_1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	out_valid;
input 	mem_used_0;
input 	mem_87_0;
input 	mem_54_0;
output 	burst_uncompress_address_base_1;
output 	burst_uncompress_address_offset_1;
input 	mem_19_0;
input 	comb;
input 	mem_57_0;
output 	source_addr_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_address_base~0_combout ;
wire \comb~0_combout ;
wire \Add2~0_combout ;
wire \p1_burst_uncompress_address_offset[0]~combout ;
wire \burst_uncompress_address_offset[0]~q ;
wire \comb~1_combout ;
wire \Add2~1 ;
wire \Add2~2_combout ;
wire \p1_burst_uncompress_address_offset[1]~combout ;


dffeas \burst_uncompress_address_base[1] (
	.clk(clk),
	.d(\burst_uncompress_address_base~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(burst_uncompress_address_base_1),
	.prn(vcc));
defparam \burst_uncompress_address_base[1] .is_wysiwyg = "true";
defparam \burst_uncompress_address_base[1] .power_up = "low";

dffeas \burst_uncompress_address_offset[1] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[1]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(burst_uncompress_address_offset_1),
	.prn(vcc));
defparam \burst_uncompress_address_offset[1] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[1] .power_up = "low";

cycloneive_lcell_comb \source_addr[1]~0 (
	.dataa(mem_19_0),
	.datab(comb),
	.datac(burst_uncompress_address_base_1),
	.datad(burst_uncompress_address_offset_1),
	.cin(gnd),
	.combout(source_addr_1),
	.cout());
defparam \source_addr[1]~0 .lut_mask = 16'hFFB8;
defparam \source_addr[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \burst_uncompress_address_base~0 (
	.dataa(mem_19_0),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_54_0),
	.cin(gnd),
	.combout(\burst_uncompress_address_base~0_combout ),
	.cout());
defparam \burst_uncompress_address_base~0 .lut_mask = 16'hAAFF;
defparam \burst_uncompress_address_base~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~0 (
	.dataa(burst_uncompress_address_offset_1),
	.datab(mem_19_0),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hAACC;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add2~0 (
	.dataa(\comb~1_combout ),
	.datab(mem_57_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
defparam \Add2~0 .lut_mask = 16'h66BB;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p1_burst_uncompress_address_offset[0] (
	.dataa(mem_54_0),
	.datab(\Add2~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p1_burst_uncompress_address_offset[0]~combout ),
	.cout());
defparam \p1_burst_uncompress_address_offset[0] .lut_mask = 16'hEEEE;
defparam \p1_burst_uncompress_address_offset[0] .sum_lutc_input = "datac";

dffeas \burst_uncompress_address_offset[0] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[0]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(\burst_uncompress_address_offset[0]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[0] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[0] .power_up = "low";

cycloneive_lcell_comb \comb~1 (
	.dataa(\burst_uncompress_address_offset[0]~q ),
	.datab(mem_87_0),
	.datac(out_valid),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(\comb~1_combout ),
	.cout());
defparam \comb~1 .lut_mask = 16'hBFFF;
defparam \comb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add2~2 (
	.dataa(\comb~0_combout ),
	.datab(mem_57_0),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout());
defparam \Add2~2 .lut_mask = 16'h9696;
defparam \Add2~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \p1_burst_uncompress_address_offset[1] (
	.dataa(mem_54_0),
	.datab(\Add2~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p1_burst_uncompress_address_offset[1]~combout ),
	.cout());
defparam \p1_burst_uncompress_address_offset[1] .lut_mask = 16'hEEEE;
defparam \p1_burst_uncompress_address_offset[1] .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_agent_11 (
	mem_used_1,
	always1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	always1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \m0_write~0 (
	.dataa(always1),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~0 .lut_mask = 16'hAAFF;
defparam \m0_write~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_agent_12 (
	mem_used_0,
	mem_105_0,
	read_latency_shift_reg_0,
	mem_used_01,
	rp_valid1,
	in_ready,
	rf_sink_ready,
	rp_valid2)/* synthesis synthesis_greybox=1 */;
input 	mem_used_0;
input 	mem_105_0;
input 	read_latency_shift_reg_0;
input 	mem_used_01;
output 	rp_valid1;
input 	in_ready;
output 	rf_sink_ready;
output 	rp_valid2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_altera_merlin_burst_uncompressor_12 uncompressor(
	.mem_used_0(mem_used_0),
	.mem_105_0(mem_105_0),
	.rp_valid(rp_valid1),
	.in_ready(in_ready),
	.sink_ready(rf_sink_ready));

cycloneive_lcell_comb \rp_valid~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(rp_valid1),
	.cout());
defparam \rp_valid~0 .lut_mask = 16'h0FFF;
defparam \rp_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb rp_valid(
	.dataa(read_latency_shift_reg_0),
	.datab(mem_used_01),
	.datac(mem_used_0),
	.datad(mem_105_0),
	.cin(gnd),
	.combout(rp_valid2),
	.cout());
defparam rp_valid.lut_mask = 16'hFFFE;
defparam rp_valid.sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_burst_uncompressor_12 (
	mem_used_0,
	mem_105_0,
	rp_valid,
	in_ready,
	sink_ready)/* synthesis synthesis_greybox=1 */;
input 	mem_used_0;
input 	mem_105_0;
input 	rp_valid;
input 	in_ready;
output 	sink_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \sink_ready~0 (
	.dataa(mem_used_0),
	.datab(mem_105_0),
	.datac(rp_valid),
	.datad(in_ready),
	.cin(gnd),
	.combout(sink_ready),
	.cout());
defparam \sink_ready~0 .lut_mask = 16'hEFFF;
defparam \sink_ready~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_agent_13 (
	hold_waitrequest,
	d_write,
	write_accepted,
	m0_write,
	Equal4,
	mem_used_1,
	m0_write1)/* synthesis synthesis_greybox=1 */;
input 	hold_waitrequest;
input 	d_write;
input 	write_accepted;
output 	m0_write;
input 	Equal4;
input 	mem_used_1;
output 	m0_write1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \m0_write~0 (
	.dataa(hold_waitrequest),
	.datab(d_write),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~0 .lut_mask = 16'hEEFF;
defparam \m0_write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_write~1 (
	.dataa(Equal4),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(m0_write1),
	.cout());
defparam \m0_write~1 .lut_mask = 16'hAAFF;
defparam \m0_write~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator (
	clk,
	reset,
	mem_used_1,
	Equal3,
	read_latency_shift_reg_0,
	always0,
	waitrequest,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_15,
	av_readdata_pre_11,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_01,
	av_readdata,
	write)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	mem_used_1;
input 	Equal3;
output 	read_latency_shift_reg_0;
input 	always0;
input 	waitrequest;
input 	read_latency_shift_reg;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_15;
output 	av_readdata_pre_11;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
output 	av_readdata_pre_01;
input 	[31:0] av_readdata;
input 	write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

cycloneive_lcell_comb \av_readdata_pre[0]~0 (
	.dataa(write),
	.datab(Equal3),
	.datac(mem_used_1),
	.datad(always0),
	.cin(gnd),
	.combout(av_readdata_pre_01),
	.cout());
defparam \av_readdata_pre[0]~0 .lut_mask = 16'hEFFF;
defparam \av_readdata_pre[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(Equal3),
	.datab(read_latency_shift_reg),
	.datac(mem_used_1),
	.datad(waitrequest),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_1 (
	clk,
	av_readdata,
	reset,
	hold_waitrequest,
	read_latency_shift_reg_0,
	write,
	mem,
	WideOr1,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_11,
	av_readdata_pre_13,
	av_readdata_pre_16,
	av_readdata_pre_12,
	av_readdata_pre_5,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_21,
	av_readdata_pre_30,
	av_readdata_pre_29,
	av_readdata_pre_28,
	av_readdata_pre_27,
	av_readdata_pre_26,
	av_readdata_pre_25,
	av_readdata_pre_24,
	av_readdata_pre_23,
	av_readdata_pre_22,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_31)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	[31:0] av_readdata;
input 	reset;
input 	hold_waitrequest;
output 	read_latency_shift_reg_0;
input 	write;
input 	mem;
input 	WideOr1;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_11;
output 	av_readdata_pre_13;
output 	av_readdata_pre_16;
output 	av_readdata_pre_12;
output 	av_readdata_pre_5;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	av_readdata_pre_21;
output 	av_readdata_pre_30;
output 	av_readdata_pre_29;
output 	av_readdata_pre_28;
output 	av_readdata_pre_27;
output 	av_readdata_pre_26;
output 	av_readdata_pre_25;
output 	av_readdata_pre_24;
output 	av_readdata_pre_23;
output 	av_readdata_pre_22;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
output 	av_readdata_pre_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(hold_waitrequest),
	.datab(write),
	.datac(WideOr1),
	.datad(mem),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_2 (
	clk,
	reset,
	wait_latency_counter_0,
	waitrequest_reset_override1,
	mem_used_1,
	wait_latency_counter_1,
	last_cycle,
	src_valid,
	src_valid1,
	p1_wr_strobe,
	src_data_66,
	av_begintransfer,
	read_latency_shift_reg_0,
	uav_waitrequest,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_11,
	av_readdata_pre_13,
	av_readdata_pre_16,
	av_readdata_pre_12,
	av_readdata_pre_5,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_21,
	av_readdata_pre_30,
	av_readdata_pre_29,
	av_readdata_pre_28,
	av_readdata_pre_27,
	av_readdata_pre_26,
	av_readdata_pre_25,
	av_readdata_pre_24,
	av_readdata_pre_23,
	av_readdata_pre_22,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata,
	av_readdata_pre_31,
	WideOr1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
output 	wait_latency_counter_0;
output 	waitrequest_reset_override1;
input 	mem_used_1;
output 	wait_latency_counter_1;
input 	last_cycle;
input 	src_valid;
input 	src_valid1;
input 	p1_wr_strobe;
input 	src_data_66;
output 	av_begintransfer;
output 	read_latency_shift_reg_0;
output 	uav_waitrequest;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_11;
output 	av_readdata_pre_13;
output 	av_readdata_pre_16;
output 	av_readdata_pre_12;
output 	av_readdata_pre_5;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	av_readdata_pre_21;
output 	av_readdata_pre_30;
output 	av_readdata_pre_29;
output 	av_readdata_pre_28;
output 	av_readdata_pre_27;
output 	av_readdata_pre_26;
output 	av_readdata_pre_25;
output 	av_readdata_pre_24;
output 	av_readdata_pre_23;
output 	av_readdata_pre_22;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
input 	[31:0] av_readdata;
output 	av_readdata_pre_31;
input 	WideOr1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas waitrequest_reset_override(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest_reset_override1),
	.prn(vcc));
defparam waitrequest_reset_override.is_wysiwyg = "true";
defparam waitrequest_reset_override.power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cycloneive_lcell_comb \av_begintransfer~0 (
	.dataa(WideOr1),
	.datab(p1_wr_strobe),
	.datac(src_data_66),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(av_begintransfer),
	.cout());
defparam \av_begintransfer~0 .lut_mask = 16'hFEFF;
defparam \av_begintransfer~0 .sum_lutc_input = "datac";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \uav_waitrequest~0 (
	.dataa(wait_latency_counter_1),
	.datab(gnd),
	.datac(wait_latency_counter_0),
	.datad(waitrequest_reset_override1),
	.cin(gnd),
	.combout(uav_waitrequest),
	.cout());
defparam \uav_waitrequest~0 .lut_mask = 16'hAFFF;
defparam \uav_waitrequest~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter~0 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(waitrequest_reset_override1),
	.datad(av_begintransfer),
	.cin(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.cout());
defparam \wait_latency_counter~0 .lut_mask = 16'hFFF5;
defparam \wait_latency_counter~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~1 (
	.dataa(wait_latency_counter_1),
	.datab(waitrequest_reset_override1),
	.datac(av_begintransfer),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.cout());
defparam \wait_latency_counter~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(last_cycle),
	.datab(src_data_66),
	.datac(src_valid),
	.datad(src_valid1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_3 (
	av_readdata_pre_22,
	av_readdata_pre_21,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_16,
	reset,
	rst1,
	b_full,
	out_data_toggle_flopped,
	av_readdata,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	dreg_0,
	av_waitrequest,
	mem_used_1,
	out_data_buffer_66,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	b_full1,
	counter_reg_bit_21,
	counter_reg_bit_11,
	counter_reg_bit_51,
	counter_reg_bit_41,
	counter_reg_bit_31,
	counter_reg_bit_01,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_15,
	av_readdata_pre_14,
	av_readdata_pre_13,
	av_readdata_pre_12,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	read_0,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_22;
output 	av_readdata_pre_21;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
output 	av_readdata_pre_16;
input 	reset;
input 	rst1;
input 	b_full;
input 	out_data_toggle_flopped;
input 	[31:0] av_readdata;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	dreg_0;
input 	av_waitrequest;
input 	mem_used_1;
input 	out_data_buffer_66;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg;
input 	b_full1;
input 	counter_reg_bit_21;
input 	counter_reg_bit_11;
input 	counter_reg_bit_51;
input 	counter_reg_bit_41;
input 	counter_reg_bit_31;
input 	counter_reg_bit_01;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_15;
output 	av_readdata_pre_14;
output 	av_readdata_pre_13;
output 	av_readdata_pre_12;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
input 	read_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \av_readdata_pre[16]~8 ;
wire \av_readdata_pre[17]~10 ;
wire \av_readdata_pre[18]~12 ;
wire \av_readdata_pre[19]~14 ;
wire \av_readdata_pre[20]~16 ;
wire \av_readdata_pre[21]~18 ;
wire \av_readdata_pre[22]~19_combout ;
wire \av_readdata_pre[21]~17_combout ;
wire \av_readdata_pre[20]~15_combout ;
wire \av_readdata_pre[19]~13_combout ;
wire \av_readdata_pre[18]~11_combout ;
wire \av_readdata_pre[17]~9_combout ;
wire \av_readdata_pre[16]~7_combout ;
wire \read_latency_shift_reg~1_combout ;
wire \av_readdata_pre[13]~21_combout ;


dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(\av_readdata_pre[22]~19_combout ),
	.asdata(b_full),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(\av_readdata_pre[21]~17_combout ),
	.asdata(counter_reg_bit_5),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(\av_readdata_pre[20]~15_combout ),
	.asdata(counter_reg_bit_4),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(\av_readdata_pre[19]~13_combout ),
	.asdata(counter_reg_bit_3),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(\av_readdata_pre[18]~11_combout ),
	.asdata(counter_reg_bit_2),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(\av_readdata_pre[17]~9_combout ),
	.asdata(counter_reg_bit_1),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(\av_readdata_pre[16]~7_combout ),
	.asdata(counter_reg_bit_0),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(av_waitrequest),
	.datab(out_data_toggle_flopped),
	.datac(dreg_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hBEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

cycloneive_lcell_comb \av_readdata_pre[16]~7 (
	.dataa(counter_reg_bit_01),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\av_readdata_pre[16]~7_combout ),
	.cout(\av_readdata_pre[16]~8 ));
defparam \av_readdata_pre[16]~7 .lut_mask = 16'hAA55;
defparam \av_readdata_pre[16]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata_pre[17]~9 (
	.dataa(counter_reg_bit_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[16]~8 ),
	.combout(\av_readdata_pre[17]~9_combout ),
	.cout(\av_readdata_pre[17]~10 ));
defparam \av_readdata_pre[17]~9 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[17]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[18]~11 (
	.dataa(counter_reg_bit_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[17]~10 ),
	.combout(\av_readdata_pre[18]~11_combout ),
	.cout(\av_readdata_pre[18]~12 ));
defparam \av_readdata_pre[18]~11 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[18]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[19]~13 (
	.dataa(counter_reg_bit_31),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[18]~12 ),
	.combout(\av_readdata_pre[19]~13_combout ),
	.cout(\av_readdata_pre[19]~14 ));
defparam \av_readdata_pre[19]~13 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[19]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[20]~15 (
	.dataa(counter_reg_bit_41),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[19]~14 ),
	.combout(\av_readdata_pre[20]~15_combout ),
	.cout(\av_readdata_pre[20]~16 ));
defparam \av_readdata_pre[20]~15 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[20]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[21]~17 (
	.dataa(counter_reg_bit_51),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[20]~16 ),
	.combout(\av_readdata_pre[21]~17_combout ),
	.cout(\av_readdata_pre[21]~18 ));
defparam \av_readdata_pre[21]~17 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[21]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[22]~19 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\av_readdata_pre[21]~18 ),
	.combout(\av_readdata_pre[22]~19_combout ),
	.cout());
defparam \av_readdata_pre[22]~19 .lut_mask = 16'h5A5A;
defparam \av_readdata_pre[22]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(rst1),
	.datab(out_data_buffer_66),
	.datac(read_latency_shift_reg),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hFEFE;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata_pre[13]~21 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_readdata_pre[13]~21_combout ),
	.cout());
defparam \av_readdata_pre[13]~21 .lut_mask = 16'h5555;
defparam \av_readdata_pre[13]~21 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_4 (
	clk,
	W_alu_result_5,
	W_alu_result_4,
	reset,
	Equal6,
	src_channel_12,
	read_latency_shift_reg_0,
	mem_used_1,
	read_latency_shift_reg,
	read_latency_shift_reg1,
	read_latency_shift_reg2)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	reset;
input 	Equal6;
input 	src_channel_12;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
output 	read_latency_shift_reg;
input 	read_latency_shift_reg1;
output 	read_latency_shift_reg2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg2),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(W_alu_result_4),
	.datab(src_channel_12),
	.datac(W_alu_result_5),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(Equal6),
	.datab(src_channel_12),
	.datac(read_latency_shift_reg1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg2),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_5 (
	clk,
	reset,
	d_read,
	read_accepted,
	hold_waitrequest,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	write)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	d_read;
input 	read_accepted;
input 	hold_waitrequest;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg;
input 	write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~3_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~2 (
	.dataa(hold_waitrequest),
	.datab(d_read),
	.datac(gnd),
	.datad(read_accepted),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~2 .lut_mask = 16'hEEFF;
defparam \read_latency_shift_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~3 (
	.dataa(hold_waitrequest),
	.datab(d_read),
	.datac(read_accepted),
	.datad(write),
	.cin(gnd),
	.combout(\read_latency_shift_reg~3_combout ),
	.cout());
defparam \read_latency_shift_reg~3 .lut_mask = 16'hFFEF;
defparam \read_latency_shift_reg~3 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_6 (
	clk,
	W_alu_result_5,
	W_alu_result_4,
	reset,
	Equal9,
	mem_used_1,
	read_latency_shift_reg,
	Equal5,
	read_latency_shift_reg_0,
	read_latency_shift_reg1,
	read_latency_shift_reg2)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	reset;
input 	Equal9;
input 	mem_used_1;
output 	read_latency_shift_reg;
input 	Equal5;
output 	read_latency_shift_reg_0;
input 	read_latency_shift_reg1;
output 	read_latency_shift_reg2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(Equal9),
	.datab(W_alu_result_5),
	.datac(W_alu_result_4),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hBFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg2),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(Equal9),
	.datab(Equal5),
	.datac(read_latency_shift_reg1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg2),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_7 (
	clk,
	reset,
	d_read,
	read_accepted,
	hold_waitrequest,
	read_latency_shift_reg_0,
	write)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	d_read;
input 	read_accepted;
input 	hold_waitrequest;
output 	read_latency_shift_reg_0;
input 	write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~2_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~2 (
	.dataa(hold_waitrequest),
	.datab(d_read),
	.datac(read_accepted),
	.datad(write),
	.cin(gnd),
	.combout(\read_latency_shift_reg~2_combout ),
	.cout());
defparam \read_latency_shift_reg~2 .lut_mask = 16'hFFEF;
defparam \read_latency_shift_reg~2 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_8 (
	clk,
	reset,
	Equal9,
	read_latency_shift_reg_0,
	mem_used_1,
	read_latency_shift_reg,
	Equal12,
	read_latency_shift_reg1,
	read_latency_shift_reg2)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	Equal9;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
input 	read_latency_shift_reg;
input 	Equal12;
output 	read_latency_shift_reg1;
output 	read_latency_shift_reg2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(Equal9),
	.datab(Equal12),
	.datac(read_latency_shift_reg),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg1),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(Equal9),
	.datab(Equal12),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg2),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hEEFF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_9 (
	clk,
	W_alu_result_3,
	reset,
	d_read,
	read_accepted,
	hold_waitrequest,
	Equal9,
	Equal6,
	read_latency_shift_reg_0,
	mem_used_1,
	read_latency_shift_reg,
	read_latency_shift_reg1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_3;
input 	reset;
input 	d_read;
input 	read_accepted;
input 	hold_waitrequest;
input 	Equal9;
input 	Equal6;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
output 	read_latency_shift_reg;
output 	read_latency_shift_reg1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~2 (
	.dataa(W_alu_result_3),
	.datab(Equal9),
	.datac(Equal6),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~2 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~3 (
	.dataa(hold_waitrequest),
	.datab(d_read),
	.datac(read_accepted),
	.datad(read_latency_shift_reg),
	.cin(gnd),
	.combout(read_latency_shift_reg1),
	.cout());
defparam \read_latency_shift_reg~3 .lut_mask = 16'hFFEF;
defparam \read_latency_shift_reg~3 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_11 (
	clk,
	W_alu_result_3,
	av_readdata,
	reset,
	uav_read,
	cp_valid,
	m0_write,
	Equal9,
	Equal6,
	read_latency_shift_reg_0,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready,
	av_waitrequest_generated,
	m0_write1,
	av_readdata_pre_30)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_3;
input 	[31:0] av_readdata;
input 	reset;
input 	uav_read;
input 	cp_valid;
input 	m0_write;
input 	Equal9;
input 	Equal6;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	sink_ready;
output 	av_waitrequest_generated;
input 	m0_write1;
output 	av_readdata_pre_30;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \av_waitrequest_generated~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cycloneive_lcell_comb \av_waitrequest_generated~1 (
	.dataa(wait_latency_counter_0),
	.datab(m0_write),
	.datac(Equal9),
	.datad(\av_waitrequest_generated~0_combout ),
	.cin(gnd),
	.combout(av_waitrequest_generated),
	.cout());
defparam \av_waitrequest_generated~1 .lut_mask = 16'h6996;
defparam \av_waitrequest_generated~1 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(cp_valid),
	.datab(m0_write1),
	.datac(wait_latency_counter_1),
	.datad(av_waitrequest_generated),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.cout());
defparam \wait_latency_counter[0]~0 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~1 (
	.dataa(\wait_latency_counter[0]~0_combout ),
	.datab(gnd),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.cout());
defparam \wait_latency_counter~1 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter[0]~0_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest_generated~0 (
	.dataa(mem_used_1),
	.datab(uav_read),
	.datac(Equal6),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\av_waitrequest_generated~0_combout ),
	.cout());
defparam \av_waitrequest_generated~0 .lut_mask = 16'hFFBF;
defparam \av_waitrequest_generated~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_12 (
	wire_pfdena_reg_ena,
	reset,
	rst1,
	out_data_buffer_66,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pfdena_reg_ena;
input 	reset;
input 	rst1;
input 	out_data_buffer_66;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(wire_pfdena_reg_ena),
	.datab(rst1),
	.datac(out_data_buffer_66),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_slave_translator_13 (
	clk,
	reset,
	cp_valid,
	m0_write,
	Equal4,
	read_latency_shift_reg_0,
	mem_used_1,
	m0_write1,
	wait_latency_counter_0,
	wait_latency_counter_1,
	read_latency_shift_reg,
	read_latency_shift_reg1,
	av_waitrequest_generated,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_15,
	av_readdata_pre_14,
	av_readdata_pre_13,
	av_readdata_pre_12,
	av_readdata_pre_11,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	cp_valid;
input 	m0_write;
input 	Equal4;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
input 	m0_write1;
output 	wait_latency_counter_0;
output 	wait_latency_counter_1;
output 	read_latency_shift_reg;
input 	read_latency_shift_reg1;
output 	av_waitrequest_generated;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_15;
output 	av_readdata_pre_14;
output 	av_readdata_pre_13;
output 	av_readdata_pre_12;
output 	av_readdata_pre_11;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
input 	[31:0] av_readdata;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~1_combout ;
wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(m0_write1),
	.datab(m0_write),
	.datac(wait_latency_counter_0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hBEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest_generated~0 (
	.dataa(wait_latency_counter_0),
	.datab(mem_used_1),
	.datac(m0_write),
	.datad(Equal4),
	.cin(gnd),
	.combout(av_waitrequest_generated),
	.cout());
defparam \av_waitrequest_generated~0 .lut_mask = 16'h6996;
defparam \av_waitrequest_generated~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(m0_write1),
	.datab(av_waitrequest_generated),
	.datac(read_latency_shift_reg1),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(cp_valid),
	.datab(m0_write1),
	.datac(wait_latency_counter_1),
	.datad(av_waitrequest_generated),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.cout());
defparam \wait_latency_counter[1]~0 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~1 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter[1]~0_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.cout());
defparam \wait_latency_counter~1 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter[1]~0_combout ),
	.datab(gnd),
	.datac(wait_latency_counter_0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_width_adapter (
	clk,
	byteen_reg_0,
	byteen_reg_1,
	address_reg_1,
	reset,
	d_writedata_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	saved_grant_0,
	use_reg1,
	WideOr0,
	Equal0,
	WideOr1,
	mem_used_7,
	src_data_46,
	out_data_28,
	src_data_60,
	out_data_42,
	src_data_47,
	out_data_29,
	src_data_49,
	out_data_31,
	src_data_48,
	out_data_30,
	src_data_51,
	out_data_33,
	src_data_50,
	out_data_32,
	src_data_53,
	out_data_35,
	src_data_52,
	out_data_34,
	src_data_55,
	out_data_37,
	src_data_54,
	out_data_36,
	src_data_57,
	out_data_39,
	src_data_56,
	out_data_38,
	src_data_59,
	out_data_41,
	src_data_58,
	out_data_40,
	out_data_19,
	src_data_38,
	out_data_20,
	src_data_39,
	out_data_21,
	src_data_40,
	out_data_22,
	src_data_41,
	out_data_23,
	src_data_42,
	out_data_24,
	src_data_43,
	out_data_25,
	src_data_44,
	out_data_26,
	src_data_45,
	out_data_27,
	count_0,
	d_writedata_10,
	in_endofpacket,
	cp_ready,
	src_data_34,
	src_data_35,
	d_writedata_8,
	d_writedata_9,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	out_endofpacket,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	byteen_reg_0;
output 	byteen_reg_1;
output 	address_reg_1;
input 	reset;
input 	d_writedata_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	saved_grant_0;
output 	use_reg1;
input 	WideOr0;
input 	Equal0;
input 	WideOr1;
input 	mem_used_7;
input 	src_data_46;
output 	out_data_28;
input 	src_data_60;
output 	out_data_42;
input 	src_data_47;
output 	out_data_29;
input 	src_data_49;
output 	out_data_31;
input 	src_data_48;
output 	out_data_30;
input 	src_data_51;
output 	out_data_33;
input 	src_data_50;
output 	out_data_32;
input 	src_data_53;
output 	out_data_35;
input 	src_data_52;
output 	out_data_34;
input 	src_data_55;
output 	out_data_37;
input 	src_data_54;
output 	out_data_36;
input 	src_data_57;
output 	out_data_39;
input 	src_data_56;
output 	out_data_38;
input 	src_data_59;
output 	out_data_41;
input 	src_data_58;
output 	out_data_40;
output 	out_data_19;
input 	src_data_38;
output 	out_data_20;
input 	src_data_39;
output 	out_data_21;
input 	src_data_40;
output 	out_data_22;
input 	src_data_41;
output 	out_data_23;
input 	src_data_42;
output 	out_data_24;
input 	src_data_43;
output 	out_data_25;
input 	src_data_44;
output 	out_data_26;
input 	src_data_45;
output 	out_data_27;
output 	count_0;
input 	d_writedata_10;
input 	in_endofpacket;
input 	cp_ready;
input 	src_data_34;
input 	src_data_35;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
output 	out_endofpacket;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_reg[11]~0_combout ;
wire \address_reg~0_combout ;
wire \use_reg~0_combout ;
wire \address_reg[10]~q ;
wire \address_reg[24]~q ;
wire \address_reg[11]~q ;
wire \address_reg[13]~q ;
wire \address_reg[12]~q ;
wire \address_reg[15]~q ;
wire \address_reg[14]~q ;
wire \address_reg[17]~q ;
wire \address_reg[16]~q ;
wire \address_reg[19]~q ;
wire \address_reg[18]~q ;
wire \address_reg[21]~q ;
wire \address_reg[20]~q ;
wire \address_reg[23]~q ;
wire \address_reg[22]~q ;
wire \address_reg[2]~q ;
wire \address_reg[3]~q ;
wire \address_reg[4]~q ;
wire \address_reg[5]~q ;
wire \address_reg[6]~q ;
wire \address_reg[7]~q ;
wire \address_reg[8]~q ;
wire \address_reg[9]~q ;
wire \count[0]~0_combout ;
wire \endofpacket_reg~q ;
wire \data_reg[0]~q ;
wire \data_reg[1]~q ;
wire \data_reg[2]~q ;
wire \data_reg[3]~q ;
wire \data_reg[4]~q ;
wire \data_reg[5]~q ;
wire \data_reg[6]~q ;
wire \data_reg[7]~q ;
wire \data_reg[8]~q ;
wire \data_reg[9]~q ;
wire \data_reg[10]~q ;
wire \data_reg[11]~q ;
wire \data_reg[12]~q ;
wire \data_reg[13]~q ;
wire \data_reg[14]~q ;
wire \data_reg[15]~q ;


dffeas \byteen_reg[0] (
	.clk(clk),
	.d(src_data_34),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(byteen_reg_0),
	.prn(vcc));
defparam \byteen_reg[0] .is_wysiwyg = "true";
defparam \byteen_reg[0] .power_up = "low";

dffeas \byteen_reg[1] (
	.clk(clk),
	.d(src_data_35),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(byteen_reg_1),
	.prn(vcc));
defparam \byteen_reg[1] .is_wysiwyg = "true";
defparam \byteen_reg[1] .power_up = "low";

dffeas \address_reg[1] (
	.clk(clk),
	.d(\address_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!use_reg1),
	.ena(vcc),
	.q(address_reg_1),
	.prn(vcc));
defparam \address_reg[1] .is_wysiwyg = "true";
defparam \address_reg[1] .power_up = "low";

dffeas use_reg(
	.clk(clk),
	.d(\use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(use_reg1),
	.prn(vcc));
defparam use_reg.is_wysiwyg = "true";
defparam use_reg.power_up = "low";

cycloneive_lcell_comb \out_data[28]~0 (
	.dataa(\address_reg[10]~q ),
	.datab(src_data_46),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_28),
	.cout());
defparam \out_data[28]~0 .lut_mask = 16'hAACC;
defparam \out_data[28]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[42]~1 (
	.dataa(\address_reg[24]~q ),
	.datab(src_data_60),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_42),
	.cout());
defparam \out_data[42]~1 .lut_mask = 16'hAACC;
defparam \out_data[42]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[29]~2 (
	.dataa(\address_reg[11]~q ),
	.datab(src_data_47),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_29),
	.cout());
defparam \out_data[29]~2 .lut_mask = 16'hAACC;
defparam \out_data[29]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[31]~3 (
	.dataa(\address_reg[13]~q ),
	.datab(src_data_49),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_31),
	.cout());
defparam \out_data[31]~3 .lut_mask = 16'hAACC;
defparam \out_data[31]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[30]~4 (
	.dataa(\address_reg[12]~q ),
	.datab(src_data_48),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_30),
	.cout());
defparam \out_data[30]~4 .lut_mask = 16'hAACC;
defparam \out_data[30]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[33]~5 (
	.dataa(\address_reg[15]~q ),
	.datab(src_data_51),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_33),
	.cout());
defparam \out_data[33]~5 .lut_mask = 16'hAACC;
defparam \out_data[33]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[32]~6 (
	.dataa(\address_reg[14]~q ),
	.datab(src_data_50),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_32),
	.cout());
defparam \out_data[32]~6 .lut_mask = 16'hAACC;
defparam \out_data[32]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[35]~7 (
	.dataa(\address_reg[17]~q ),
	.datab(src_data_53),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_35),
	.cout());
defparam \out_data[35]~7 .lut_mask = 16'hAACC;
defparam \out_data[35]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[34]~8 (
	.dataa(\address_reg[16]~q ),
	.datab(src_data_52),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_34),
	.cout());
defparam \out_data[34]~8 .lut_mask = 16'hAACC;
defparam \out_data[34]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[37]~9 (
	.dataa(\address_reg[19]~q ),
	.datab(src_data_55),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_37),
	.cout());
defparam \out_data[37]~9 .lut_mask = 16'hAACC;
defparam \out_data[37]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[36]~10 (
	.dataa(\address_reg[18]~q ),
	.datab(src_data_54),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_36),
	.cout());
defparam \out_data[36]~10 .lut_mask = 16'hAACC;
defparam \out_data[36]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[39]~11 (
	.dataa(\address_reg[21]~q ),
	.datab(src_data_57),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_39),
	.cout());
defparam \out_data[39]~11 .lut_mask = 16'hAACC;
defparam \out_data[39]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[38]~12 (
	.dataa(\address_reg[20]~q ),
	.datab(src_data_56),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_38),
	.cout());
defparam \out_data[38]~12 .lut_mask = 16'hAACC;
defparam \out_data[38]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[41]~13 (
	.dataa(\address_reg[23]~q ),
	.datab(src_data_59),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_41),
	.cout());
defparam \out_data[41]~13 .lut_mask = 16'hAACC;
defparam \out_data[41]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[40]~14 (
	.dataa(\address_reg[22]~q ),
	.datab(src_data_58),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_40),
	.cout());
defparam \out_data[40]~14 .lut_mask = 16'hAACC;
defparam \out_data[40]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[19]~15 (
	.dataa(use_reg1),
	.datab(address_reg_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_data_19),
	.cout());
defparam \out_data[19]~15 .lut_mask = 16'hEEEE;
defparam \out_data[19]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[20]~16 (
	.dataa(\address_reg[2]~q ),
	.datab(src_data_38),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_20),
	.cout());
defparam \out_data[20]~16 .lut_mask = 16'hAACC;
defparam \out_data[20]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[21]~17 (
	.dataa(\address_reg[3]~q ),
	.datab(src_data_39),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_21),
	.cout());
defparam \out_data[21]~17 .lut_mask = 16'hAACC;
defparam \out_data[21]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[22]~18 (
	.dataa(\address_reg[4]~q ),
	.datab(src_data_40),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_22),
	.cout());
defparam \out_data[22]~18 .lut_mask = 16'hAACC;
defparam \out_data[22]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[23]~19 (
	.dataa(\address_reg[5]~q ),
	.datab(src_data_41),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_23),
	.cout());
defparam \out_data[23]~19 .lut_mask = 16'hAACC;
defparam \out_data[23]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[24]~20 (
	.dataa(\address_reg[6]~q ),
	.datab(src_data_42),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_24),
	.cout());
defparam \out_data[24]~20 .lut_mask = 16'hAACC;
defparam \out_data[24]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[25]~21 (
	.dataa(\address_reg[7]~q ),
	.datab(src_data_43),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_25),
	.cout());
defparam \out_data[25]~21 .lut_mask = 16'hAACC;
defparam \out_data[25]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[26]~22 (
	.dataa(\address_reg[8]~q ),
	.datab(src_data_44),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_26),
	.cout());
defparam \out_data[26]~22 .lut_mask = 16'hAACC;
defparam \out_data[26]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[27]~23 (
	.dataa(\address_reg[9]~q ),
	.datab(src_data_45),
	.datac(gnd),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_27),
	.cout());
defparam \out_data[27]~23 .lut_mask = 16'hAACC;
defparam \out_data[27]~23 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(count_0),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneive_lcell_comb \out_endofpacket~0 (
	.dataa(use_reg1),
	.datab(count_0),
	.datac(\endofpacket_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(out_endofpacket),
	.cout());
defparam \out_endofpacket~0 .lut_mask = 16'hFEFE;
defparam \out_endofpacket~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[0]~24 (
	.dataa(\data_reg[0]~q ),
	.datab(d_writedata_0),
	.datac(saved_grant_0),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_0),
	.cout());
defparam \out_data[0]~24 .lut_mask = 16'hFAFC;
defparam \out_data[0]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[1]~25 (
	.dataa(\data_reg[1]~q ),
	.datab(d_writedata_1),
	.datac(saved_grant_0),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_1),
	.cout());
defparam \out_data[1]~25 .lut_mask = 16'hFAFC;
defparam \out_data[1]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[2]~26 (
	.dataa(\data_reg[2]~q ),
	.datab(d_writedata_2),
	.datac(saved_grant_0),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_2),
	.cout());
defparam \out_data[2]~26 .lut_mask = 16'hFAFC;
defparam \out_data[2]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[3]~27 (
	.dataa(\data_reg[3]~q ),
	.datab(d_writedata_3),
	.datac(saved_grant_0),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_3),
	.cout());
defparam \out_data[3]~27 .lut_mask = 16'hFAFC;
defparam \out_data[3]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[4]~28 (
	.dataa(\data_reg[4]~q ),
	.datab(d_writedata_4),
	.datac(saved_grant_0),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_4),
	.cout());
defparam \out_data[4]~28 .lut_mask = 16'hFAFC;
defparam \out_data[4]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[5]~29 (
	.dataa(\data_reg[5]~q ),
	.datab(d_writedata_5),
	.datac(saved_grant_0),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_5),
	.cout());
defparam \out_data[5]~29 .lut_mask = 16'hFAFC;
defparam \out_data[5]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[6]~30 (
	.dataa(\data_reg[6]~q ),
	.datab(d_writedata_6),
	.datac(saved_grant_0),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_6),
	.cout());
defparam \out_data[6]~30 .lut_mask = 16'hFAFC;
defparam \out_data[6]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[7]~31 (
	.dataa(\data_reg[7]~q ),
	.datab(d_writedata_7),
	.datac(saved_grant_0),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_7),
	.cout());
defparam \out_data[7]~31 .lut_mask = 16'hFAFC;
defparam \out_data[7]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[8]~32 (
	.dataa(\data_reg[8]~q ),
	.datab(saved_grant_0),
	.datac(d_writedata_8),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_8),
	.cout());
defparam \out_data[8]~32 .lut_mask = 16'hFAFC;
defparam \out_data[8]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[9]~33 (
	.dataa(\data_reg[9]~q ),
	.datab(saved_grant_0),
	.datac(d_writedata_9),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_9),
	.cout());
defparam \out_data[9]~33 .lut_mask = 16'hFAFC;
defparam \out_data[9]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[10]~34 (
	.dataa(\data_reg[10]~q ),
	.datab(saved_grant_0),
	.datac(d_writedata_10),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_10),
	.cout());
defparam \out_data[10]~34 .lut_mask = 16'hFAFC;
defparam \out_data[10]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[11]~35 (
	.dataa(\data_reg[11]~q ),
	.datab(saved_grant_0),
	.datac(d_writedata_11),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_11),
	.cout());
defparam \out_data[11]~35 .lut_mask = 16'hFAFC;
defparam \out_data[11]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[12]~36 (
	.dataa(\data_reg[12]~q ),
	.datab(saved_grant_0),
	.datac(d_writedata_12),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_12),
	.cout());
defparam \out_data[12]~36 .lut_mask = 16'hFAFC;
defparam \out_data[12]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[13]~37 (
	.dataa(\data_reg[13]~q ),
	.datab(saved_grant_0),
	.datac(d_writedata_13),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_13),
	.cout());
defparam \out_data[13]~37 .lut_mask = 16'hFAFC;
defparam \out_data[13]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[14]~38 (
	.dataa(\data_reg[14]~q ),
	.datab(saved_grant_0),
	.datac(d_writedata_14),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_14),
	.cout());
defparam \out_data[14]~38 .lut_mask = 16'hFAFC;
defparam \out_data[14]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[15]~39 (
	.dataa(\data_reg[15]~q ),
	.datab(saved_grant_0),
	.datac(d_writedata_15),
	.datad(use_reg1),
	.cin(gnd),
	.combout(out_data_15),
	.cout());
defparam \out_data[15]~39 .lut_mask = 16'hFAFC;
defparam \out_data[15]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg[11]~0 (
	.dataa(use_reg1),
	.datab(mem_used_7),
	.datac(Equal0),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\data_reg[11]~0_combout ),
	.cout());
defparam \data_reg[11]~0 .lut_mask = 16'h7FFF;
defparam \data_reg[11]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_reg~0 (
	.dataa(Equal0),
	.datab(WideOr0),
	.datac(mem_used_7),
	.datad(address_reg_1),
	.cin(gnd),
	.combout(\address_reg~0_combout ),
	.cout());
defparam \address_reg~0 .lut_mask = 16'h6996;
defparam \address_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \use_reg~0 (
	.dataa(use_reg1),
	.datab(cp_ready),
	.datac(WideOr1),
	.datad(count_0),
	.cin(gnd),
	.combout(\use_reg~0_combout ),
	.cout());
defparam \use_reg~0 .lut_mask = 16'hF6FF;
defparam \use_reg~0 .sum_lutc_input = "datac";

dffeas \address_reg[10] (
	.clk(clk),
	.d(src_data_46),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[10]~q ),
	.prn(vcc));
defparam \address_reg[10] .is_wysiwyg = "true";
defparam \address_reg[10] .power_up = "low";

dffeas \address_reg[24] (
	.clk(clk),
	.d(src_data_60),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[24]~q ),
	.prn(vcc));
defparam \address_reg[24] .is_wysiwyg = "true";
defparam \address_reg[24] .power_up = "low";

dffeas \address_reg[11] (
	.clk(clk),
	.d(src_data_47),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[11]~q ),
	.prn(vcc));
defparam \address_reg[11] .is_wysiwyg = "true";
defparam \address_reg[11] .power_up = "low";

dffeas \address_reg[13] (
	.clk(clk),
	.d(src_data_49),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[13]~q ),
	.prn(vcc));
defparam \address_reg[13] .is_wysiwyg = "true";
defparam \address_reg[13] .power_up = "low";

dffeas \address_reg[12] (
	.clk(clk),
	.d(src_data_48),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[12]~q ),
	.prn(vcc));
defparam \address_reg[12] .is_wysiwyg = "true";
defparam \address_reg[12] .power_up = "low";

dffeas \address_reg[15] (
	.clk(clk),
	.d(src_data_51),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[15]~q ),
	.prn(vcc));
defparam \address_reg[15] .is_wysiwyg = "true";
defparam \address_reg[15] .power_up = "low";

dffeas \address_reg[14] (
	.clk(clk),
	.d(src_data_50),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[14]~q ),
	.prn(vcc));
defparam \address_reg[14] .is_wysiwyg = "true";
defparam \address_reg[14] .power_up = "low";

dffeas \address_reg[17] (
	.clk(clk),
	.d(src_data_53),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[17]~q ),
	.prn(vcc));
defparam \address_reg[17] .is_wysiwyg = "true";
defparam \address_reg[17] .power_up = "low";

dffeas \address_reg[16] (
	.clk(clk),
	.d(src_data_52),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[16]~q ),
	.prn(vcc));
defparam \address_reg[16] .is_wysiwyg = "true";
defparam \address_reg[16] .power_up = "low";

dffeas \address_reg[19] (
	.clk(clk),
	.d(src_data_55),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[19]~q ),
	.prn(vcc));
defparam \address_reg[19] .is_wysiwyg = "true";
defparam \address_reg[19] .power_up = "low";

dffeas \address_reg[18] (
	.clk(clk),
	.d(src_data_54),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[18]~q ),
	.prn(vcc));
defparam \address_reg[18] .is_wysiwyg = "true";
defparam \address_reg[18] .power_up = "low";

dffeas \address_reg[21] (
	.clk(clk),
	.d(src_data_57),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[21]~q ),
	.prn(vcc));
defparam \address_reg[21] .is_wysiwyg = "true";
defparam \address_reg[21] .power_up = "low";

dffeas \address_reg[20] (
	.clk(clk),
	.d(src_data_56),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[20]~q ),
	.prn(vcc));
defparam \address_reg[20] .is_wysiwyg = "true";
defparam \address_reg[20] .power_up = "low";

dffeas \address_reg[23] (
	.clk(clk),
	.d(src_data_59),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[23]~q ),
	.prn(vcc));
defparam \address_reg[23] .is_wysiwyg = "true";
defparam \address_reg[23] .power_up = "low";

dffeas \address_reg[22] (
	.clk(clk),
	.d(src_data_58),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[22]~q ),
	.prn(vcc));
defparam \address_reg[22] .is_wysiwyg = "true";
defparam \address_reg[22] .power_up = "low";

dffeas \address_reg[2] (
	.clk(clk),
	.d(src_data_38),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[2]~q ),
	.prn(vcc));
defparam \address_reg[2] .is_wysiwyg = "true";
defparam \address_reg[2] .power_up = "low";

dffeas \address_reg[3] (
	.clk(clk),
	.d(src_data_39),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[3]~q ),
	.prn(vcc));
defparam \address_reg[3] .is_wysiwyg = "true";
defparam \address_reg[3] .power_up = "low";

dffeas \address_reg[4] (
	.clk(clk),
	.d(src_data_40),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[4]~q ),
	.prn(vcc));
defparam \address_reg[4] .is_wysiwyg = "true";
defparam \address_reg[4] .power_up = "low";

dffeas \address_reg[5] (
	.clk(clk),
	.d(src_data_41),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[5]~q ),
	.prn(vcc));
defparam \address_reg[5] .is_wysiwyg = "true";
defparam \address_reg[5] .power_up = "low";

dffeas \address_reg[6] (
	.clk(clk),
	.d(src_data_42),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[6]~q ),
	.prn(vcc));
defparam \address_reg[6] .is_wysiwyg = "true";
defparam \address_reg[6] .power_up = "low";

dffeas \address_reg[7] (
	.clk(clk),
	.d(src_data_43),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[7]~q ),
	.prn(vcc));
defparam \address_reg[7] .is_wysiwyg = "true";
defparam \address_reg[7] .power_up = "low";

dffeas \address_reg[8] (
	.clk(clk),
	.d(src_data_44),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[8]~q ),
	.prn(vcc));
defparam \address_reg[8] .is_wysiwyg = "true";
defparam \address_reg[8] .power_up = "low";

dffeas \address_reg[9] (
	.clk(clk),
	.d(src_data_45),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\address_reg[9]~q ),
	.prn(vcc));
defparam \address_reg[9] .is_wysiwyg = "true";
defparam \address_reg[9] .power_up = "low";

cycloneive_lcell_comb \count[0]~0 (
	.dataa(count_0),
	.datab(cp_ready),
	.datac(WideOr1),
	.datad(use_reg1),
	.cin(gnd),
	.combout(\count[0]~0_combout ),
	.cout());
defparam \count[0]~0 .lut_mask = 16'hF9F6;
defparam \count[0]~0 .sum_lutc_input = "datac";

dffeas endofpacket_reg(
	.clk(clk),
	.d(in_endofpacket),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!use_reg1),
	.q(\endofpacket_reg~q ),
	.prn(vcc));
defparam endofpacket_reg.is_wysiwyg = "true";
defparam endofpacket_reg.power_up = "low";

dffeas \data_reg[0] (
	.clk(clk),
	.d(src_payload),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[0]~q ),
	.prn(vcc));
defparam \data_reg[0] .is_wysiwyg = "true";
defparam \data_reg[0] .power_up = "low";

dffeas \data_reg[1] (
	.clk(clk),
	.d(src_payload1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[1]~q ),
	.prn(vcc));
defparam \data_reg[1] .is_wysiwyg = "true";
defparam \data_reg[1] .power_up = "low";

dffeas \data_reg[2] (
	.clk(clk),
	.d(src_payload2),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[2]~q ),
	.prn(vcc));
defparam \data_reg[2] .is_wysiwyg = "true";
defparam \data_reg[2] .power_up = "low";

dffeas \data_reg[3] (
	.clk(clk),
	.d(src_payload3),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[3]~q ),
	.prn(vcc));
defparam \data_reg[3] .is_wysiwyg = "true";
defparam \data_reg[3] .power_up = "low";

dffeas \data_reg[4] (
	.clk(clk),
	.d(src_payload4),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[4]~q ),
	.prn(vcc));
defparam \data_reg[4] .is_wysiwyg = "true";
defparam \data_reg[4] .power_up = "low";

dffeas \data_reg[5] (
	.clk(clk),
	.d(src_payload5),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[5]~q ),
	.prn(vcc));
defparam \data_reg[5] .is_wysiwyg = "true";
defparam \data_reg[5] .power_up = "low";

dffeas \data_reg[6] (
	.clk(clk),
	.d(src_payload6),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[6]~q ),
	.prn(vcc));
defparam \data_reg[6] .is_wysiwyg = "true";
defparam \data_reg[6] .power_up = "low";

dffeas \data_reg[7] (
	.clk(clk),
	.d(src_payload7),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[7]~q ),
	.prn(vcc));
defparam \data_reg[7] .is_wysiwyg = "true";
defparam \data_reg[7] .power_up = "low";

dffeas \data_reg[8] (
	.clk(clk),
	.d(src_payload8),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[8]~q ),
	.prn(vcc));
defparam \data_reg[8] .is_wysiwyg = "true";
defparam \data_reg[8] .power_up = "low";

dffeas \data_reg[9] (
	.clk(clk),
	.d(src_payload9),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[9]~q ),
	.prn(vcc));
defparam \data_reg[9] .is_wysiwyg = "true";
defparam \data_reg[9] .power_up = "low";

dffeas \data_reg[10] (
	.clk(clk),
	.d(src_payload10),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[10]~q ),
	.prn(vcc));
defparam \data_reg[10] .is_wysiwyg = "true";
defparam \data_reg[10] .power_up = "low";

dffeas \data_reg[11] (
	.clk(clk),
	.d(src_payload11),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[11]~q ),
	.prn(vcc));
defparam \data_reg[11] .is_wysiwyg = "true";
defparam \data_reg[11] .power_up = "low";

dffeas \data_reg[12] (
	.clk(clk),
	.d(src_payload12),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[12]~q ),
	.prn(vcc));
defparam \data_reg[12] .is_wysiwyg = "true";
defparam \data_reg[12] .power_up = "low";

dffeas \data_reg[13] (
	.clk(clk),
	.d(src_payload13),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[13]~q ),
	.prn(vcc));
defparam \data_reg[13] .is_wysiwyg = "true";
defparam \data_reg[13] .power_up = "low";

dffeas \data_reg[14] (
	.clk(clk),
	.d(src_payload14),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[14]~q ),
	.prn(vcc));
defparam \data_reg[14] .is_wysiwyg = "true";
defparam \data_reg[14] .power_up = "low";

dffeas \data_reg[15] (
	.clk(clk),
	.d(src_payload15),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(use_reg1),
	.sload(gnd),
	.ena(\data_reg[11]~0_combout ),
	.q(\data_reg[15]~q ),
	.prn(vcc));
defparam \data_reg[15] .is_wysiwyg = "true";
defparam \data_reg[15] .power_up = "low";

endmodule

module niosII_altera_merlin_width_adapter_1 (
	wire_pll7_clk_0,
	r_sync_rst,
	rp_valid,
	mem_88_0,
	mem_54_0,
	burst_uncompress_address_base_1,
	burst_uncompress_address_offset_1,
	mem_19_0,
	comb,
	always10,
	data_reg_0,
	out_payload_0,
	source_addr_1,
	data_reg_1,
	out_payload_1,
	data_reg_2,
	out_payload_2,
	data_reg_3,
	out_payload_3,
	data_reg_4,
	out_payload_4,
	data_reg_11,
	out_payload_11,
	data_reg_13,
	out_payload_13,
	data_reg_12,
	out_payload_12,
	data_reg_5,
	out_payload_5,
	data_reg_14,
	out_payload_14,
	data_reg_15,
	out_payload_15,
	data_reg_10,
	out_payload_10,
	data_reg_9,
	out_payload_9,
	data_reg_8,
	out_payload_8,
	data_reg_7,
	out_payload_7,
	data_reg_6,
	out_payload_6)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	rp_valid;
input 	mem_88_0;
input 	mem_54_0;
input 	burst_uncompress_address_base_1;
input 	burst_uncompress_address_offset_1;
input 	mem_19_0;
input 	comb;
output 	always10;
output 	data_reg_0;
input 	out_payload_0;
input 	source_addr_1;
output 	data_reg_1;
input 	out_payload_1;
output 	data_reg_2;
input 	out_payload_2;
output 	data_reg_3;
input 	out_payload_3;
output 	data_reg_4;
input 	out_payload_4;
output 	data_reg_11;
input 	out_payload_11;
output 	data_reg_13;
input 	out_payload_13;
output 	data_reg_12;
input 	out_payload_12;
output 	data_reg_5;
input 	out_payload_5;
output 	data_reg_14;
input 	out_payload_14;
output 	data_reg_15;
input 	out_payload_15;
output 	data_reg_10;
input 	out_payload_10;
output 	data_reg_9;
input 	out_payload_9;
output 	data_reg_8;
input 	out_payload_8;
output 	data_reg_7;
input 	out_payload_7;
output 	data_reg_6;
input 	out_payload_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always10~0_combout ;
wire \data_reg~0_combout ;
wire \data_reg~1_combout ;
wire \data_reg~2_combout ;
wire \data_reg~3_combout ;
wire \data_reg~4_combout ;
wire \data_reg~5_combout ;
wire \data_reg~6_combout ;
wire \data_reg~7_combout ;
wire \data_reg~8_combout ;
wire \data_reg~9_combout ;
wire \data_reg~10_combout ;
wire \data_reg~11_combout ;
wire \data_reg~12_combout ;
wire \data_reg~13_combout ;
wire \data_reg~14_combout ;
wire \data_reg~15_combout ;


cycloneive_lcell_comb \always10~1 (
	.dataa(mem_88_0),
	.datab(mem_54_0),
	.datac(\always10~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(always10),
	.cout());
defparam \always10~1 .lut_mask = 16'hFBFB;
defparam \always10~1 .sum_lutc_input = "datac";

dffeas \data_reg[0] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_0),
	.prn(vcc));
defparam \data_reg[0] .is_wysiwyg = "true";
defparam \data_reg[0] .power_up = "low";

dffeas \data_reg[1] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_1),
	.prn(vcc));
defparam \data_reg[1] .is_wysiwyg = "true";
defparam \data_reg[1] .power_up = "low";

dffeas \data_reg[2] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_2),
	.prn(vcc));
defparam \data_reg[2] .is_wysiwyg = "true";
defparam \data_reg[2] .power_up = "low";

dffeas \data_reg[3] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_3),
	.prn(vcc));
defparam \data_reg[3] .is_wysiwyg = "true";
defparam \data_reg[3] .power_up = "low";

dffeas \data_reg[4] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_4),
	.prn(vcc));
defparam \data_reg[4] .is_wysiwyg = "true";
defparam \data_reg[4] .power_up = "low";

dffeas \data_reg[11] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_11),
	.prn(vcc));
defparam \data_reg[11] .is_wysiwyg = "true";
defparam \data_reg[11] .power_up = "low";

dffeas \data_reg[13] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_13),
	.prn(vcc));
defparam \data_reg[13] .is_wysiwyg = "true";
defparam \data_reg[13] .power_up = "low";

dffeas \data_reg[12] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_12),
	.prn(vcc));
defparam \data_reg[12] .is_wysiwyg = "true";
defparam \data_reg[12] .power_up = "low";

dffeas \data_reg[5] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_5),
	.prn(vcc));
defparam \data_reg[5] .is_wysiwyg = "true";
defparam \data_reg[5] .power_up = "low";

dffeas \data_reg[14] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_14),
	.prn(vcc));
defparam \data_reg[14] .is_wysiwyg = "true";
defparam \data_reg[14] .power_up = "low";

dffeas \data_reg[15] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_15),
	.prn(vcc));
defparam \data_reg[15] .is_wysiwyg = "true";
defparam \data_reg[15] .power_up = "low";

dffeas \data_reg[10] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_10),
	.prn(vcc));
defparam \data_reg[10] .is_wysiwyg = "true";
defparam \data_reg[10] .power_up = "low";

dffeas \data_reg[9] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_9),
	.prn(vcc));
defparam \data_reg[9] .is_wysiwyg = "true";
defparam \data_reg[9] .power_up = "low";

dffeas \data_reg[8] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_8),
	.prn(vcc));
defparam \data_reg[8] .is_wysiwyg = "true";
defparam \data_reg[8] .power_up = "low";

dffeas \data_reg[7] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_7),
	.prn(vcc));
defparam \data_reg[7] .is_wysiwyg = "true";
defparam \data_reg[7] .power_up = "low";

dffeas \data_reg[6] (
	.clk(wire_pll7_clk_0),
	.d(\data_reg~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rp_valid),
	.q(data_reg_6),
	.prn(vcc));
defparam \data_reg[6] .is_wysiwyg = "true";
defparam \data_reg[6] .power_up = "low";

cycloneive_lcell_comb \always10~0 (
	.dataa(burst_uncompress_address_base_1),
	.datab(burst_uncompress_address_offset_1),
	.datac(mem_19_0),
	.datad(comb),
	.cin(gnd),
	.combout(\always10~0_combout ),
	.cout());
defparam \always10~0 .lut_mask = 16'hFAFC;
defparam \always10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~0 (
	.dataa(data_reg_0),
	.datab(out_payload_0),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~0_combout ),
	.cout());
defparam \data_reg~0 .lut_mask = 16'hEFFF;
defparam \data_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~1 (
	.dataa(data_reg_1),
	.datab(out_payload_1),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~1_combout ),
	.cout());
defparam \data_reg~1 .lut_mask = 16'hEFFF;
defparam \data_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~2 (
	.dataa(data_reg_2),
	.datab(out_payload_2),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~2_combout ),
	.cout());
defparam \data_reg~2 .lut_mask = 16'hEFFF;
defparam \data_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~3 (
	.dataa(data_reg_3),
	.datab(out_payload_3),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~3_combout ),
	.cout());
defparam \data_reg~3 .lut_mask = 16'hEFFF;
defparam \data_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~4 (
	.dataa(data_reg_4),
	.datab(out_payload_4),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~4_combout ),
	.cout());
defparam \data_reg~4 .lut_mask = 16'hEFFF;
defparam \data_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~5 (
	.dataa(data_reg_11),
	.datab(out_payload_11),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~5_combout ),
	.cout());
defparam \data_reg~5 .lut_mask = 16'hEFFF;
defparam \data_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~6 (
	.dataa(data_reg_13),
	.datab(out_payload_13),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~6_combout ),
	.cout());
defparam \data_reg~6 .lut_mask = 16'hEFFF;
defparam \data_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~7 (
	.dataa(data_reg_12),
	.datab(out_payload_12),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~7_combout ),
	.cout());
defparam \data_reg~7 .lut_mask = 16'hEFFF;
defparam \data_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~8 (
	.dataa(data_reg_5),
	.datab(out_payload_5),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~8_combout ),
	.cout());
defparam \data_reg~8 .lut_mask = 16'hEFFF;
defparam \data_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~9 (
	.dataa(data_reg_14),
	.datab(out_payload_14),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~9_combout ),
	.cout());
defparam \data_reg~9 .lut_mask = 16'hEFFF;
defparam \data_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~10 (
	.dataa(data_reg_15),
	.datab(out_payload_15),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~10_combout ),
	.cout());
defparam \data_reg~10 .lut_mask = 16'hEFFF;
defparam \data_reg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~11 (
	.dataa(data_reg_10),
	.datab(out_payload_10),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~11_combout ),
	.cout());
defparam \data_reg~11 .lut_mask = 16'hEFFF;
defparam \data_reg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~12 (
	.dataa(data_reg_9),
	.datab(out_payload_9),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~12_combout ),
	.cout());
defparam \data_reg~12 .lut_mask = 16'hEFFF;
defparam \data_reg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~13 (
	.dataa(data_reg_8),
	.datab(out_payload_8),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~13_combout ),
	.cout());
defparam \data_reg~13 .lut_mask = 16'hEFFF;
defparam \data_reg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~14 (
	.dataa(data_reg_7),
	.datab(out_payload_7),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~14_combout ),
	.cout());
defparam \data_reg~14 .lut_mask = 16'hEFFF;
defparam \data_reg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~15 (
	.dataa(data_reg_6),
	.datab(out_payload_6),
	.datac(source_addr_1),
	.datad(always10),
	.cin(gnd),
	.combout(\data_reg~15_combout ),
	.cout());
defparam \data_reg~15 .lut_mask = 16'hEFFF;
defparam \data_reg~15 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_mm_interconnect_0_cmd_demux (
	W_alu_result_5,
	W_alu_result_4,
	hold_waitrequest,
	d_write,
	write_accepted,
	cp_valid,
	Equal9,
	mem_used_1,
	saved_grant_0,
	src_channel_12,
	Equal2,
	src_channel_121,
	src_channel_122,
	Equal1,
	src_channel_123,
	src12_valid,
	waitrequest,
	m0_read,
	last_cycle,
	in_ready,
	src_channel_124,
	WideOr0,
	read_latency_shift_reg,
	read_latency_shift_reg1,
	mem_used_11,
	mem_used_12,
	write,
	Equal12,
	mem_used_13,
	mem_used_14,
	wait_latency_counter_1,
	always1,
	wait_latency_counter_0,
	sink_ready,
	take_in_data,
	saved_grant_01,
	waitrequest1,
	mem_used_15,
	Equal13,
	in_data_toggle,
	dreg_0,
	WideOr01,
	src12_valid1,
	av_waitrequest_generated,
	sink_ready1)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	hold_waitrequest;
input 	d_write;
input 	write_accepted;
input 	cp_valid;
input 	Equal9;
input 	mem_used_1;
input 	saved_grant_0;
input 	src_channel_12;
input 	Equal2;
input 	src_channel_121;
input 	src_channel_122;
input 	Equal1;
input 	src_channel_123;
output 	src12_valid;
input 	waitrequest;
input 	m0_read;
input 	last_cycle;
input 	in_ready;
input 	src_channel_124;
output 	WideOr0;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg1;
input 	mem_used_11;
input 	mem_used_12;
input 	write;
input 	Equal12;
input 	mem_used_13;
input 	mem_used_14;
input 	wait_latency_counter_1;
input 	always1;
input 	wait_latency_counter_0;
output 	sink_ready;
input 	take_in_data;
input 	saved_grant_01;
input 	waitrequest1;
input 	mem_used_15;
input 	Equal13;
input 	in_data_toggle;
input 	dreg_0;
output 	WideOr01;
output 	src12_valid1;
input 	av_waitrequest_generated;
output 	sink_ready1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~0_combout ;
wire \sink_ready~5_combout ;
wire \WideOr0~2_combout ;
wire \WideOr0~3_combout ;
wire \WideOr0~4_combout ;
wire \WideOr0~5_combout ;
wire \WideOr0~6_combout ;
wire \sink_ready~3_combout ;
wire \WideOr0~7_combout ;
wire \src12_valid~1_combout ;


cycloneive_lcell_comb \src12_valid~0 (
	.dataa(cp_valid),
	.datab(src_channel_12),
	.datac(src_channel_123),
	.datad(src_channel_122),
	.cin(gnd),
	.combout(src12_valid),
	.cout());
defparam \src12_valid~0 .lut_mask = 16'hBFFF;
defparam \src12_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~1 (
	.dataa(m0_read),
	.datab(\WideOr0~0_combout ),
	.datac(waitrequest),
	.datad(src_channel_124),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hEFFF;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~2 (
	.dataa(mem_used_14),
	.datab(wait_latency_counter_1),
	.datac(always1),
	.datad(\sink_ready~5_combout ),
	.cin(gnd),
	.combout(sink_ready),
	.cout());
defparam \sink_ready~2 .lut_mask = 16'hFFF7;
defparam \sink_ready~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~8 (
	.dataa(\WideOr0~6_combout ),
	.datab(sink_ready),
	.datac(take_in_data),
	.datad(\WideOr0~7_combout ),
	.cin(gnd),
	.combout(WideOr01),
	.cout());
defparam \WideOr0~8 .lut_mask = 16'hFFFE;
defparam \WideOr0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src12_valid~2 (
	.dataa(src_channel_12),
	.datab(src_channel_123),
	.datac(src_channel_122),
	.datad(\src12_valid~1_combout ),
	.cin(gnd),
	.combout(src12_valid1),
	.cout());
defparam \src12_valid~2 .lut_mask = 16'hFF7F;
defparam \src12_valid~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~4 (
	.dataa(hold_waitrequest),
	.datab(always1),
	.datac(av_waitrequest_generated),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(sink_ready1),
	.cout());
defparam \sink_ready~4 .lut_mask = 16'hFEFF;
defparam \sink_ready~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(saved_grant_0),
	.datab(last_cycle),
	.datac(Equal1),
	.datad(in_ready),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hACFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~5 (
	.dataa(hold_waitrequest),
	.datab(d_write),
	.datac(write_accepted),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\sink_ready~5_combout ),
	.cout());
defparam \sink_ready~5 .lut_mask = 16'hEBBE;
defparam \sink_ready~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~2 (
	.dataa(mem_used_11),
	.datab(W_alu_result_5),
	.datac(W_alu_result_4),
	.datad(mem_used_12),
	.cin(gnd),
	.combout(\WideOr0~2_combout ),
	.cout());
defparam \WideOr0~2 .lut_mask = 16'h7DFF;
defparam \WideOr0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~3 (
	.dataa(W_alu_result_4),
	.datab(mem_used_1),
	.datac(\WideOr0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr0~3_combout ),
	.cout());
defparam \WideOr0~3 .lut_mask = 16'hFBFB;
defparam \WideOr0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~4 (
	.dataa(Equal9),
	.datab(W_alu_result_4),
	.datac(src_channel_121),
	.datad(\WideOr0~3_combout ),
	.cin(gnd),
	.combout(\WideOr0~4_combout ),
	.cout());
defparam \WideOr0~4 .lut_mask = 16'hFFB8;
defparam \WideOr0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~5 (
	.dataa(\WideOr0~4_combout ),
	.datab(write),
	.datac(Equal12),
	.datad(mem_used_13),
	.cin(gnd),
	.combout(\WideOr0~5_combout ),
	.cout());
defparam \WideOr0~5 .lut_mask = 16'hFEFF;
defparam \WideOr0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~6 (
	.dataa(hold_waitrequest),
	.datab(read_latency_shift_reg),
	.datac(read_latency_shift_reg1),
	.datad(\WideOr0~5_combout ),
	.cin(gnd),
	.combout(\WideOr0~6_combout ),
	.cout());
defparam \WideOr0~6 .lut_mask = 16'hFFFE;
defparam \WideOr0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~3 (
	.dataa(Equal2),
	.datab(saved_grant_01),
	.datac(waitrequest1),
	.datad(mem_used_15),
	.cin(gnd),
	.combout(\sink_ready~3_combout ),
	.cout());
defparam \sink_ready~3 .lut_mask = 16'hEFFF;
defparam \sink_ready~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~7 (
	.dataa(\sink_ready~3_combout ),
	.datab(Equal13),
	.datac(in_data_toggle),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\WideOr0~7_combout ),
	.cout());
defparam \WideOr0~7 .lut_mask = 16'hEFFE;
defparam \WideOr0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src12_valid~1 (
	.dataa(cp_valid),
	.datab(Equal1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src12_valid~1_combout ),
	.cout());
defparam \src12_valid~1 .lut_mask = 16'hBBBB;
defparam \src12_valid~1 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_mm_interconnect_0_cmd_demux_001 (
	hold_waitrequest,
	i_read,
	read_accepted,
	Equal1,
	uav_read,
	F_pc_9,
	src0_valid,
	src2_valid)/* synthesis synthesis_greybox=1 */;
input 	hold_waitrequest;
input 	i_read;
input 	read_accepted;
input 	Equal1;
input 	uav_read;
input 	F_pc_9;
output 	src0_valid;
output 	src2_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(hold_waitrequest),
	.datab(uav_read),
	.datac(F_pc_9),
	.datad(Equal1),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hFFFE;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src2_valid~2 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(hold_waitrequest),
	.datad(Equal1),
	.cin(gnd),
	.combout(src2_valid),
	.cout());
defparam \src2_valid~2 .lut_mask = 16'hF7FF;
defparam \src2_valid~2 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_mm_interconnect_0_cmd_mux_009 (
	wire_pll7_clk_0,
	W_alu_result_6,
	W_alu_result_10,
	W_alu_result_5,
	W_alu_result_7,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	r_sync_rst,
	cp_valid,
	d_writedata_0,
	d_byteenable_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_byteenable_1,
	Equal2,
	F_pc_8,
	F_pc_0,
	F_pc_1,
	F_pc_2,
	F_pc_3,
	F_pc_4,
	F_pc_5,
	F_pc_6,
	F_pc_7,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	d_writedata_10,
	d_byteenable_2,
	d_byteenable_3,
	saved_grant_1,
	hbreak_enabled,
	d_writedata_8,
	d_writedata_9,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	src0_valid,
	WideOr11,
	src_data_46,
	src_payload,
	src_payload1,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_data_33,
	src_payload7,
	src_payload8,
	src_data_34,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_data_35,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_6;
input 	W_alu_result_10;
input 	W_alu_result_5;
input 	W_alu_result_7;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	r_sync_rst;
input 	cp_valid;
input 	d_writedata_0;
input 	d_byteenable_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_byteenable_1;
input 	Equal2;
input 	F_pc_8;
input 	F_pc_0;
input 	F_pc_1;
input 	F_pc_2;
input 	F_pc_3;
input 	F_pc_4;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_7;
output 	saved_grant_0;
input 	waitrequest;
input 	mem_used_1;
input 	d_writedata_10;
input 	d_byteenable_2;
input 	d_byteenable_3;
output 	saved_grant_1;
input 	hbreak_enabled;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
input 	src0_valid;
output 	WideOr11;
output 	src_data_46;
output 	src_payload;
output 	src_payload1;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_32;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_data_33;
output 	src_payload7;
output 	src_payload8;
output 	src_data_34;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_data_35;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~0_combout ;


niosII_altera_merlin_arbitrator arb(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.cp_valid(cp_valid),
	.Equal2(Equal2),
	.src0_valid(src0_valid),
	.src_valid(\src_valid~0_combout ),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ));

dffeas \saved_grant[0] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(src0_valid),
	.datad(\src_valid~0_combout ),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[46] (
	.dataa(W_alu_result_10),
	.datab(F_pc_8),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(d_writedata_0),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[40] (
	.dataa(W_alu_result_4),
	.datab(F_pc_2),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[41] (
	.dataa(W_alu_result_5),
	.datab(F_pc_3),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[42] (
	.dataa(W_alu_result_6),
	.datab(F_pc_4),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[43] (
	.dataa(W_alu_result_7),
	.datab(F_pc_5),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[44] (
	.dataa(W_alu_result_8),
	.datab(F_pc_6),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[45] (
	.dataa(W_alu_result_9),
	.datab(F_pc_7),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[32] (
	.dataa(saved_grant_1),
	.datab(d_byteenable_0),
	.datac(saved_grant_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_32),
	.cout());
defparam \src_data[32] .lut_mask = 16'hFEFE;
defparam \src_data[32] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(d_writedata_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(d_writedata_4),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(d_writedata_3),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(d_writedata_2),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(saved_grant_0),
	.datab(d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[33] (
	.dataa(saved_grant_1),
	.datab(d_byteenable_1),
	.datac(saved_grant_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_33),
	.cout());
defparam \src_data[33] .lut_mask = 16'hFEFE;
defparam \src_data[33] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(saved_grant_0),
	.datab(d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[34] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_2),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_34),
	.cout());
defparam \src_data[34] .lut_mask = 16'hFEFE;
defparam \src_data[34] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(d_writedata_5),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(saved_grant_0),
	.datab(d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(saved_grant_0),
	.datab(d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(d_writedata_7),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(d_writedata_6),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(saved_grant_0),
	.datab(d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(saved_grant_0),
	.datab(d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[35] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_3),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_35),
	.cout());
defparam \src_data[35] .lut_mask = 16'hFEFE;
defparam \src_data[35] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(saved_grant_0),
	.datab(d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~21 (
	.dataa(saved_grant_0),
	.datab(d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~22 (
	.dataa(saved_grant_0),
	.datab(d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~23 (
	.dataa(saved_grant_0),
	.datab(d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~24 (
	.dataa(saved_grant_0),
	.datab(d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~25 (
	.dataa(saved_grant_0),
	.datab(d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~26 (
	.dataa(saved_grant_0),
	.datab(d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~27 (
	.dataa(saved_grant_0),
	.datab(d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~28 (
	.dataa(saved_grant_0),
	.datab(d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~29 (
	.dataa(saved_grant_0),
	.datab(d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~30 (
	.dataa(saved_grant_0),
	.datab(d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~32 (
	.dataa(saved_grant_0),
	.datab(d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload32),
	.cout());
defparam \src_payload~32 .lut_mask = 16'hEEEE;
defparam \src_payload~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEFFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(wire_pll7_clk_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(gnd),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h88BB;
defparam \update_grant~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(cp_valid),
	.datab(Equal2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~0_combout ),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hEEEE;
defparam \src_valid~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_arbitrator (
	clk,
	reset,
	cp_valid,
	Equal2,
	src0_valid,
	src_valid,
	grant_0,
	update_grant,
	grant_1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	cp_valid;
input 	Equal2;
input 	src0_valid;
input 	src_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~3_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src0_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(src0_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(\top_priority_reg[0]~q ),
	.datad(src_valid),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~2 (
	.dataa(cp_valid),
	.datab(Equal2),
	.datac(update_grant),
	.datad(src0_valid),
	.cin(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.cout());
defparam \top_priority_reg[0]~2 .lut_mask = 16'hFFFE;
defparam \top_priority_reg[0]~2 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~2_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~3 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~3_combout ),
	.cout());
defparam \top_priority_reg[0]~3 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~3 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~2_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module niosII_niosII_mm_interconnect_0_cmd_mux_009_1 (
	wire_pll7_clk_0,
	r_sync_rst,
	saved_grant_0,
	saved_grant_1,
	out_data_buffer_38,
	out_data_buffer_381,
	src_data_38,
	out_data_buffer_39,
	out_data_buffer_391,
	src_data_39,
	out_data_buffer_40,
	out_data_buffer_401,
	src_data_40,
	out_data_buffer_10,
	src_payload,
	out_data_buffer_0,
	src_payload1,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	out_data_toggle_flopped1,
	dreg_01,
	out_valid1,
	wait_latency_counter_0,
	waitrequest_reset_override,
	mem_used_1,
	wait_latency_counter_1,
	last_cycle,
	out_data_buffer_105,
	out_data_buffer_1051,
	src_payload_0,
	src_valid,
	src_valid1,
	out_data_buffer_46,
	out_data_buffer_461,
	src_data_46,
	out_data_buffer_7,
	src_payload2,
	src_payload3,
	out_data_buffer_66,
	out_data_buffer_661,
	src_data_66,
	out_data_buffer_6,
	src_payload4,
	out_data_buffer_5,
	src_payload5,
	out_data_buffer_4,
	src_payload6,
	out_data_buffer_3,
	src_payload7,
	out_data_buffer_2,
	src_payload8,
	out_data_buffer_1,
	src_payload9,
	out_data_buffer_41,
	out_data_buffer_411,
	src_data_41,
	out_data_buffer_42,
	out_data_buffer_421,
	src_data_42,
	out_data_buffer_43,
	out_data_buffer_431,
	src_data_43,
	out_data_buffer_44,
	out_data_buffer_441,
	src_data_44,
	out_data_buffer_45,
	out_data_buffer_451,
	src_data_45,
	src_payload10,
	out_data_buffer_11,
	src_payload11,
	out_data_buffer_13,
	src_payload12,
	out_data_buffer_12,
	src_payload13,
	out_data_buffer_14,
	src_payload14,
	out_data_buffer_15,
	src_payload15,
	out_data_buffer_9,
	src_payload16,
	out_data_buffer_8,
	src_payload17,
	WideOr11)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
output 	saved_grant_0;
output 	saved_grant_1;
input 	out_data_buffer_38;
input 	out_data_buffer_381;
output 	src_data_38;
input 	out_data_buffer_39;
input 	out_data_buffer_391;
output 	src_data_39;
input 	out_data_buffer_40;
input 	out_data_buffer_401;
output 	src_data_40;
input 	out_data_buffer_10;
output 	src_payload;
input 	out_data_buffer_0;
output 	src_payload1;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid;
input 	out_data_toggle_flopped1;
input 	dreg_01;
input 	out_valid1;
input 	wait_latency_counter_0;
input 	waitrequest_reset_override;
input 	mem_used_1;
input 	wait_latency_counter_1;
output 	last_cycle;
input 	out_data_buffer_105;
input 	out_data_buffer_1051;
output 	src_payload_0;
output 	src_valid;
output 	src_valid1;
input 	out_data_buffer_46;
input 	out_data_buffer_461;
output 	src_data_46;
input 	out_data_buffer_7;
output 	src_payload2;
output 	src_payload3;
input 	out_data_buffer_66;
input 	out_data_buffer_661;
output 	src_data_66;
input 	out_data_buffer_6;
output 	src_payload4;
input 	out_data_buffer_5;
output 	src_payload5;
input 	out_data_buffer_4;
output 	src_payload6;
input 	out_data_buffer_3;
output 	src_payload7;
input 	out_data_buffer_2;
output 	src_payload8;
input 	out_data_buffer_1;
output 	src_payload9;
input 	out_data_buffer_41;
input 	out_data_buffer_411;
output 	src_data_41;
input 	out_data_buffer_42;
input 	out_data_buffer_421;
output 	src_data_42;
input 	out_data_buffer_43;
input 	out_data_buffer_431;
output 	src_data_43;
input 	out_data_buffer_44;
input 	out_data_buffer_441;
output 	src_data_44;
input 	out_data_buffer_45;
input 	out_data_buffer_451;
output 	src_data_45;
output 	src_payload10;
input 	out_data_buffer_11;
output 	src_payload11;
input 	out_data_buffer_13;
output 	src_payload12;
input 	out_data_buffer_12;
output 	src_payload13;
input 	out_data_buffer_14;
output 	src_payload14;
input 	out_data_buffer_15;
output 	src_payload15;
input 	out_data_buffer_9;
output 	src_payload16;
input 	out_data_buffer_8;
output 	src_payload17;
output 	WideOr11;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


niosII_altera_merlin_arbitrator_1 arb(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.out_data_toggle_flopped(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid(out_valid),
	.out_valid1(out_valid1),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~0_combout ),
	.grant_1(\arb|grant[1]~1_combout ));

dffeas \saved_grant[0] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb \src_data[38] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_38),
	.datad(out_data_buffer_381),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_39),
	.datad(out_data_buffer_391),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[40] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_40),
	.datad(out_data_buffer_401),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \last_cycle~0 (
	.dataa(wait_latency_counter_0),
	.datab(waitrequest_reset_override),
	.datac(mem_used_1),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(last_cycle),
	.cout());
defparam \last_cycle~0 .lut_mask = 16'hEFFF;
defparam \last_cycle~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_105),
	.datad(out_data_buffer_1051),
	.cin(gnd),
	.combout(src_payload_0),
	.cout());
defparam \src_payload[0] .lut_mask = 16'hFFFE;
defparam \src_payload[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(saved_grant_0),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hAFFA;
defparam \src_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~1 (
	.dataa(saved_grant_1),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_01),
	.cin(gnd),
	.combout(src_valid1),
	.cout());
defparam \src_valid~1 .lut_mask = 16'hAFFA;
defparam \src_valid~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[46] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_46),
	.datad(out_data_buffer_461),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_381),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[66] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_66),
	.datad(out_data_buffer_661),
	.cin(gnd),
	.combout(src_data_66),
	.cout());
defparam \src_data[66] .lut_mask = 16'hFFFE;
defparam \src_data[66] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[41] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_41),
	.datad(out_data_buffer_411),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[42] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_42),
	.datad(out_data_buffer_421),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[43] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_43),
	.datad(out_data_buffer_431),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[44] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_44),
	.datad(out_data_buffer_441),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[45] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_45),
	.datad(out_data_buffer_451),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(saved_grant_1),
	.datab(out_data_buffer_38),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_0),
	.datab(out_data_toggle_flopped),
	.datac(dreg_0),
	.datad(src_valid1),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFBE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(wire_pll7_clk_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(last_cycle),
	.datab(src_payload_0),
	.datac(WideOr11),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hACFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_arbitrator_1 (
	clk,
	reset,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	out_valid1,
	grant_0,
	update_grant,
	grant_1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid;
input 	out_valid1;
output 	grant_0;
input 	update_grant;
output 	grant_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~4_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~5_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(out_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(out_valid1),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(out_valid1),
	.datab(\top_priority_reg[1]~q ),
	.datac(out_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~4 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(update_grant),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\top_priority_reg[0]~4_combout ),
	.cout());
defparam \top_priority_reg[0]~4 .lut_mask = 16'hFFF6;
defparam \top_priority_reg[0]~4 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~4_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~5 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~5_combout ),
	.cout());
defparam \top_priority_reg[0]~5 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~5 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~4_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module niosII_niosII_mm_interconnect_0_cmd_mux_009_2 (
	wire_pll7_clk_0,
	W_alu_result_6,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_5,
	W_alu_result_7,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	r_sync_rst,
	uav_read,
	cp_valid,
	saved_grant_0,
	saved_grant_1,
	WideOr0,
	Equal0,
	src_channel_12,
	src_channel_121,
	cp_valid1,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	Equal1,
	Equal11,
	src_channel_122,
	WideOr11,
	mem_used_7,
	uav_read1,
	src_data_66,
	F_pc_8,
	src_data_46,
	src_valid,
	src_data_60,
	F_pc_9,
	src_data_47,
	src_data_49,
	src_data_48,
	src_data_51,
	src_data_50,
	src_data_53,
	src_data_52,
	src_data_55,
	src_data_54,
	src_data_57,
	src_data_56,
	src_data_59,
	src_data_58,
	F_pc_0,
	src_data_38,
	F_pc_1,
	src_data_39,
	F_pc_2,
	src_data_40,
	F_pc_3,
	src_data_41,
	F_pc_4,
	src_data_42,
	F_pc_5,
	src_data_43,
	F_pc_6,
	src_data_44,
	F_pc_7,
	src_data_45,
	count_0,
	last_cycle,
	src12_valid,
	src_payload_0,
	d_byteenable_2,
	src_data_34,
	d_byteenable_3,
	src_data_35,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src2_valid)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_6;
input 	W_alu_result_24;
input 	W_alu_result_23;
input 	W_alu_result_22;
input 	W_alu_result_21;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_5;
input 	W_alu_result_7;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	r_sync_rst;
input 	uav_read;
input 	cp_valid;
output 	saved_grant_0;
output 	saved_grant_1;
input 	WideOr0;
input 	Equal0;
input 	src_channel_12;
input 	src_channel_121;
input 	cp_valid1;
input 	F_pc_22;
input 	F_pc_21;
input 	F_pc_20;
input 	F_pc_19;
input 	F_pc_18;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
input 	F_pc_10;
input 	Equal1;
input 	Equal11;
input 	src_channel_122;
output 	WideOr11;
input 	mem_used_7;
input 	uav_read1;
output 	src_data_66;
input 	F_pc_8;
output 	src_data_46;
output 	src_valid;
output 	src_data_60;
input 	F_pc_9;
output 	src_data_47;
output 	src_data_49;
output 	src_data_48;
output 	src_data_51;
output 	src_data_50;
output 	src_data_53;
output 	src_data_52;
output 	src_data_55;
output 	src_data_54;
output 	src_data_57;
output 	src_data_56;
output 	src_data_59;
output 	src_data_58;
input 	F_pc_0;
output 	src_data_38;
input 	F_pc_1;
output 	src_data_39;
input 	F_pc_2;
output 	src_data_40;
input 	F_pc_3;
output 	src_data_41;
input 	F_pc_4;
output 	src_data_42;
input 	F_pc_5;
output 	src_data_43;
input 	F_pc_6;
output 	src_data_44;
input 	F_pc_7;
output 	src_data_45;
input 	count_0;
output 	last_cycle;
input 	src12_valid;
output 	src_payload_0;
input 	d_byteenable_2;
output 	src_data_34;
input 	d_byteenable_3;
output 	src_data_35;
input 	d_writedata_16;
input 	d_writedata_17;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
input 	src2_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \WideOr1~0_combout ;
wire \WideOr1~1_combout ;


niosII_altera_merlin_arbitrator_2 arb(
	.clk(wire_pll7_clk_0),
	.reset(r_sync_rst),
	.src12_valid(src12_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~0_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src2_valid(src2_valid));

dffeas \saved_grant[0] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(src_channel_12),
	.datab(src_channel_121),
	.datac(\WideOr1~0_combout ),
	.datad(\WideOr1~1_combout ),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFF7;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[66] (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_66),
	.cout());
defparam \src_data[66] .lut_mask = 16'hFFFE;
defparam \src_data[66] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[46] (
	.dataa(W_alu_result_10),
	.datab(saved_grant_1),
	.datac(F_pc_8),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(saved_grant_1),
	.datab(cp_valid1),
	.datac(gnd),
	.datad(Equal1),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hEEFF;
defparam \src_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[60] (
	.dataa(W_alu_result_24),
	.datab(saved_grant_1),
	.datac(F_pc_22),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_60),
	.cout());
defparam \src_data[60] .lut_mask = 16'hFFFE;
defparam \src_data[60] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[47] (
	.dataa(W_alu_result_11),
	.datab(saved_grant_1),
	.datac(F_pc_9),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_47),
	.cout());
defparam \src_data[47] .lut_mask = 16'hFFFE;
defparam \src_data[47] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[49] (
	.dataa(W_alu_result_13),
	.datab(saved_grant_1),
	.datac(F_pc_11),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_49),
	.cout());
defparam \src_data[49] .lut_mask = 16'hFFFE;
defparam \src_data[49] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[48] (
	.dataa(W_alu_result_12),
	.datab(saved_grant_0),
	.datac(saved_grant_1),
	.datad(F_pc_10),
	.cin(gnd),
	.combout(src_data_48),
	.cout());
defparam \src_data[48] .lut_mask = 16'hFEFF;
defparam \src_data[48] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[51] (
	.dataa(W_alu_result_15),
	.datab(saved_grant_1),
	.datac(F_pc_13),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_51),
	.cout());
defparam \src_data[51] .lut_mask = 16'hFFFE;
defparam \src_data[51] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[50] (
	.dataa(W_alu_result_14),
	.datab(saved_grant_1),
	.datac(F_pc_12),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_50),
	.cout());
defparam \src_data[50] .lut_mask = 16'hFFFE;
defparam \src_data[50] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[53] (
	.dataa(W_alu_result_17),
	.datab(saved_grant_1),
	.datac(F_pc_15),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_53),
	.cout());
defparam \src_data[53] .lut_mask = 16'hFFFE;
defparam \src_data[53] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[52] (
	.dataa(W_alu_result_16),
	.datab(saved_grant_1),
	.datac(F_pc_14),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_52),
	.cout());
defparam \src_data[52] .lut_mask = 16'hFFFE;
defparam \src_data[52] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[55] (
	.dataa(W_alu_result_19),
	.datab(saved_grant_1),
	.datac(F_pc_17),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_55),
	.cout());
defparam \src_data[55] .lut_mask = 16'hFFFE;
defparam \src_data[55] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[54] (
	.dataa(W_alu_result_18),
	.datab(saved_grant_1),
	.datac(F_pc_16),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_54),
	.cout());
defparam \src_data[54] .lut_mask = 16'hFFFE;
defparam \src_data[54] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[57] (
	.dataa(W_alu_result_21),
	.datab(saved_grant_1),
	.datac(F_pc_19),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_57),
	.cout());
defparam \src_data[57] .lut_mask = 16'hFFFE;
defparam \src_data[57] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[56] (
	.dataa(W_alu_result_20),
	.datab(saved_grant_1),
	.datac(F_pc_18),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_56),
	.cout());
defparam \src_data[56] .lut_mask = 16'hFFFE;
defparam \src_data[56] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[59] (
	.dataa(W_alu_result_23),
	.datab(saved_grant_1),
	.datac(F_pc_21),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_59),
	.cout());
defparam \src_data[59] .lut_mask = 16'hFFFE;
defparam \src_data[59] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[58] (
	.dataa(W_alu_result_22),
	.datab(saved_grant_1),
	.datac(F_pc_20),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_58),
	.cout());
defparam \src_data[58] .lut_mask = 16'hFFFE;
defparam \src_data[58] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(saved_grant_1),
	.datac(F_pc_0),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(saved_grant_1),
	.datac(F_pc_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[40] (
	.dataa(W_alu_result_4),
	.datab(saved_grant_1),
	.datac(F_pc_2),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[41] (
	.dataa(W_alu_result_5),
	.datab(saved_grant_1),
	.datac(F_pc_3),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[42] (
	.dataa(W_alu_result_6),
	.datab(saved_grant_1),
	.datac(F_pc_4),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[43] (
	.dataa(W_alu_result_7),
	.datab(saved_grant_1),
	.datac(F_pc_5),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[44] (
	.dataa(W_alu_result_8),
	.datab(saved_grant_1),
	.datac(F_pc_6),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[45] (
	.dataa(W_alu_result_9),
	.datab(saved_grant_1),
	.datac(F_pc_7),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cycloneive_lcell_comb \last_cycle~0 (
	.dataa(count_0),
	.datab(Equal0),
	.datac(WideOr0),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(last_cycle),
	.cout());
defparam \last_cycle~0 .lut_mask = 16'hBFFF;
defparam \last_cycle~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload_0),
	.cout());
defparam \src_payload[0] .lut_mask = 16'hEEEE;
defparam \src_payload[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[34] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_2),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_34),
	.cout());
defparam \src_data[34] .lut_mask = 16'hFEFE;
defparam \src_data[34] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[35] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_3),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_35),
	.cout());
defparam \src_data[35] .lut_mask = 16'hFEFE;
defparam \src_data[35] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(saved_grant_0),
	.datab(d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(saved_grant_0),
	.datab(d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(saved_grant_0),
	.datab(d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(saved_grant_0),
	.datab(d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(saved_grant_0),
	.datab(d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(saved_grant_0),
	.datab(d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(saved_grant_0),
	.datab(d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(saved_grant_0),
	.datab(d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(saved_grant_0),
	.datab(d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(saved_grant_0),
	.datab(d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(wire_pll7_clk_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(last_cycle),
	.datab(src_payload_0),
	.datac(WideOr11),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hACFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~0 (
	.dataa(saved_grant_1),
	.datab(cp_valid1),
	.datac(Equal1),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hEFEF;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~1 (
	.dataa(saved_grant_0),
	.datab(Equal11),
	.datac(cp_valid),
	.datad(src_channel_122),
	.cin(gnd),
	.combout(\WideOr1~1_combout ),
	.cout());
defparam \WideOr1~1 .lut_mask = 16'hFBFF;
defparam \WideOr1~1 .sum_lutc_input = "datac";

endmodule

module niosII_altera_merlin_arbitrator_2 (
	clk,
	reset,
	src12_valid,
	grant_0,
	update_grant,
	grant_1,
	src2_valid)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	src12_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	src2_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(src12_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src2_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(src2_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src12_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src12_valid),
	.datac(src2_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module niosII_niosII_mm_interconnect_0_router (
	W_alu_result_6,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_5,
	W_alu_result_7,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_4,
	W_alu_result_3,
	uav_read,
	Equal3,
	Equal9,
	Equal6,
	src_channel_12,
	Equal2,
	src_channel_121,
	src_channel_122,
	Equal1,
	Equal4,
	Equal5,
	src_channel_123,
	src_channel_124,
	Equal12,
	always1,
	Equal13,
	Equal121,
	Equal51)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_6;
input 	W_alu_result_26;
input 	W_alu_result_25;
input 	W_alu_result_24;
input 	W_alu_result_23;
input 	W_alu_result_22;
input 	W_alu_result_21;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_5;
input 	W_alu_result_7;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	uav_read;
output 	Equal3;
output 	Equal9;
output 	Equal6;
output 	src_channel_12;
output 	Equal2;
output 	src_channel_121;
output 	src_channel_122;
output 	Equal1;
output 	Equal4;
output 	Equal5;
output 	src_channel_123;
output 	src_channel_124;
output 	Equal12;
output 	always1;
output 	Equal13;
output 	Equal121;
output 	Equal51;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal3~0_combout ;
wire \Equal3~1_combout ;
wire \Equal3~2_combout ;
wire \Equal3~3_combout ;
wire \Equal3~4_combout ;
wire \Equal3~5_combout ;
wire \Equal3~7_combout ;
wire \Equal2~0_combout ;
wire \src_channel[12]~2_combout ;
wire \Equal4~0_combout ;
wire \Equal12~0_combout ;
wire \Equal13~0_combout ;
wire \Equal5~1_combout ;


cycloneive_lcell_comb \Equal3~6 (
	.dataa(W_alu_result_6),
	.datab(\Equal3~3_combout ),
	.datac(\Equal3~4_combout ),
	.datad(\Equal3~5_combout ),
	.cin(gnd),
	.combout(Equal3),
	.cout());
defparam \Equal3~6 .lut_mask = 16'hFFFD;
defparam \Equal3~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal9~0 (
	.dataa(W_alu_result_7),
	.datab(\Equal3~3_combout ),
	.datac(\Equal3~7_combout ),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(Equal9),
	.cout());
defparam \Equal9~0 .lut_mask = 16'hFEFF;
defparam \Equal9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~0 (
	.dataa(W_alu_result_4),
	.datab(gnd),
	.datac(gnd),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(Equal6),
	.cout());
defparam \Equal6~0 .lut_mask = 16'hAAFF;
defparam \Equal6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[12]~0 (
	.dataa(Equal9),
	.datab(Equal6),
	.datac(uav_read),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(src_channel_12),
	.cout());
defparam \src_channel[12]~0 .lut_mask = 16'hFFFE;
defparam \src_channel[12]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~1 (
	.dataa(\Equal3~0_combout ),
	.datab(\Equal3~1_combout ),
	.datac(\Equal3~2_combout ),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hFFFE;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[12]~1 (
	.dataa(W_alu_result_6),
	.datab(\Equal3~3_combout ),
	.datac(\Equal3~7_combout ),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(src_channel_121),
	.cout());
defparam \src_channel[12]~1 .lut_mask = 16'hFEFF;
defparam \src_channel[12]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[12]~3 (
	.dataa(Equal9),
	.datab(Equal2),
	.datac(src_channel_121),
	.datad(\src_channel[12]~2_combout ),
	.cin(gnd),
	.combout(src_channel_122),
	.cout());
defparam \src_channel[12]~3 .lut_mask = 16'hFFFE;
defparam \src_channel[12]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\Equal3~3_combout ),
	.datab(W_alu_result_12),
	.datac(W_alu_result_13),
	.datad(W_alu_result_11),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal4~1 (
	.dataa(W_alu_result_5),
	.datab(\Equal3~3_combout ),
	.datac(\Equal3~4_combout ),
	.datad(\Equal4~0_combout ),
	.cin(gnd),
	.combout(Equal4),
	.cout());
defparam \Equal4~1 .lut_mask = 16'hFFFE;
defparam \Equal4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(W_alu_result_5),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(Equal5),
	.cout());
defparam \Equal5~0 .lut_mask = 16'h0FFF;
defparam \Equal5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[12]~4 (
	.dataa(Equal3),
	.datab(Equal4),
	.datac(Equal9),
	.datad(Equal5),
	.cin(gnd),
	.combout(src_channel_123),
	.cout());
defparam \src_channel[12]~4 .lut_mask = 16'hFFFE;
defparam \src_channel[12]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[12]~5 (
	.dataa(src_channel_12),
	.datab(src_channel_123),
	.datac(src_channel_122),
	.datad(gnd),
	.cin(gnd),
	.combout(src_channel_124),
	.cout());
defparam \src_channel[12]~5 .lut_mask = 16'hFEFE;
defparam \src_channel[12]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal12~1 (
	.dataa(W_alu_result_5),
	.datab(\Equal3~3_combout ),
	.datac(\Equal3~7_combout ),
	.datad(\Equal12~0_combout ),
	.cin(gnd),
	.combout(Equal12),
	.cout());
defparam \Equal12~1 .lut_mask = 16'hFFFE;
defparam \Equal12~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(uav_read),
	.datab(Equal9),
	.datac(Equal6),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(always1),
	.cout());
defparam \always1~0 .lut_mask = 16'hFEFF;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal13~1 (
	.dataa(W_alu_result_3),
	.datab(\Equal3~3_combout ),
	.datac(\Equal3~7_combout ),
	.datad(\Equal13~0_combout ),
	.cin(gnd),
	.combout(Equal13),
	.cout());
defparam \Equal13~1 .lut_mask = 16'hFFFE;
defparam \Equal13~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal12~2 (
	.dataa(W_alu_result_5),
	.datab(gnd),
	.datac(W_alu_result_4),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(Equal121),
	.cout());
defparam \Equal12~2 .lut_mask = 16'hAFFF;
defparam \Equal12~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~2 (
	.dataa(W_alu_result_5),
	.datab(\Equal3~3_combout ),
	.datac(\Equal3~7_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(Equal51),
	.cout());
defparam \Equal5~2 .lut_mask = 16'hFFFD;
defparam \Equal5~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~0 (
	.dataa(W_alu_result_26),
	.datab(W_alu_result_25),
	.datac(W_alu_result_24),
	.datad(W_alu_result_23),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
defparam \Equal3~0 .lut_mask = 16'hBFFF;
defparam \Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~1 (
	.dataa(W_alu_result_22),
	.datab(W_alu_result_21),
	.datac(W_alu_result_20),
	.datad(W_alu_result_19),
	.cin(gnd),
	.combout(\Equal3~1_combout ),
	.cout());
defparam \Equal3~1 .lut_mask = 16'h7FFF;
defparam \Equal3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~2 (
	.dataa(W_alu_result_18),
	.datab(W_alu_result_17),
	.datac(W_alu_result_16),
	.datad(W_alu_result_15),
	.cin(gnd),
	.combout(\Equal3~2_combout ),
	.cout());
defparam \Equal3~2 .lut_mask = 16'h7FFF;
defparam \Equal3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~3 (
	.dataa(\Equal3~0_combout ),
	.datab(\Equal3~1_combout ),
	.datac(\Equal3~2_combout ),
	.datad(W_alu_result_14),
	.cin(gnd),
	.combout(\Equal3~3_combout ),
	.cout());
defparam \Equal3~3 .lut_mask = 16'hFEFF;
defparam \Equal3~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~4 (
	.dataa(W_alu_result_13),
	.datab(W_alu_result_12),
	.datac(W_alu_result_11),
	.datad(W_alu_result_10),
	.cin(gnd),
	.combout(\Equal3~4_combout ),
	.cout());
defparam \Equal3~4 .lut_mask = 16'hBFFF;
defparam \Equal3~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~5 (
	.dataa(W_alu_result_5),
	.datab(W_alu_result_7),
	.datac(W_alu_result_9),
	.datad(W_alu_result_8),
	.cin(gnd),
	.combout(\Equal3~5_combout ),
	.cout());
defparam \Equal3~5 .lut_mask = 16'h7FFF;
defparam \Equal3~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~7 (
	.dataa(\Equal3~4_combout ),
	.datab(gnd),
	.datac(W_alu_result_9),
	.datad(W_alu_result_8),
	.cin(gnd),
	.combout(\Equal3~7_combout ),
	.cout());
defparam \Equal3~7 .lut_mask = 16'hAFFF;
defparam \Equal3~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(W_alu_result_12),
	.datab(W_alu_result_11),
	.datac(W_alu_result_13),
	.datad(W_alu_result_14),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hEFFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[12]~2 (
	.dataa(W_alu_result_5),
	.datab(W_alu_result_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_channel[12]~2_combout ),
	.cout());
defparam \src_channel[12]~2 .lut_mask = 16'hBBBB;
defparam \src_channel[12]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal4~0 (
	.dataa(W_alu_result_7),
	.datab(W_alu_result_6),
	.datac(W_alu_result_9),
	.datad(W_alu_result_8),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'h7FFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal12~0 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_3),
	.datac(W_alu_result_7),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(\Equal12~0_combout ),
	.cout());
defparam \Equal12~0 .lut_mask = 16'hF7FF;
defparam \Equal12~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal13~0 (
	.dataa(W_alu_result_5),
	.datab(W_alu_result_4),
	.datac(W_alu_result_7),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(\Equal13~0_combout ),
	.cout());
defparam \Equal13~0 .lut_mask = 16'hFBFF;
defparam \Equal13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~1 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_6),
	.datac(W_alu_result_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal5~1_combout ),
	.cout());
defparam \Equal5~1 .lut_mask = 16'hDFDF;
defparam \Equal5~1 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_mm_interconnect_0_router_001 (
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	Equal1)/* synthesis synthesis_greybox=1 */;
input 	F_pc_24;
input 	F_pc_23;
input 	F_pc_22;
input 	F_pc_21;
input 	F_pc_20;
input 	F_pc_19;
input 	F_pc_18;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
input 	F_pc_10;
output 	Equal1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \Equal1~2_combout ;
wire \Equal1~3_combout ;


cycloneive_lcell_comb \Equal1~4 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\Equal1~2_combout ),
	.datad(\Equal1~3_combout ),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~4 .lut_mask = 16'hFFFE;
defparam \Equal1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(F_pc_24),
	.datab(F_pc_23),
	.datac(F_pc_22),
	.datad(F_pc_21),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h7FFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(F_pc_20),
	.datab(F_pc_19),
	.datac(F_pc_18),
	.datad(F_pc_17),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'h7FFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(F_pc_16),
	.datab(F_pc_15),
	.datac(F_pc_14),
	.datad(F_pc_13),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'h7FFF;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~3 (
	.dataa(gnd),
	.datab(F_pc_12),
	.datac(F_pc_11),
	.datad(F_pc_10),
	.cin(gnd),
	.combout(\Equal1~3_combout ),
	.cout());
defparam \Equal1~3 .lut_mask = 16'h3FFF;
defparam \Equal1~3 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_mm_interconnect_0_rsp_demux_009 (
	mem_84_0,
	mem_66_0,
	read_latency_shift_reg_0,
	src1_valid,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	mem_84_0;
input 	mem_66_0;
input 	read_latency_shift_reg_0;
output 	src1_valid;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_84_0),
	.datac(mem_66_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_mm_interconnect_0_rsp_demux_009_1 (
	mem_84_0,
	mem_66_0,
	in_data_toggle,
	dreg_0,
	in_data_toggle1,
	dreg_01,
	take_in_data,
	WideOr0)/* synthesis synthesis_greybox=1 */;
input 	mem_84_0;
input 	mem_66_0;
input 	in_data_toggle;
input 	dreg_0;
input 	in_data_toggle1;
input 	dreg_01;
input 	take_in_data;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~0_combout ;


cycloneive_lcell_comb \WideOr0~1 (
	.dataa(\WideOr0~0_combout ),
	.datab(in_data_toggle1),
	.datac(dreg_01),
	.datad(take_in_data),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hBEFF;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(mem_84_0),
	.datab(mem_66_0),
	.datac(in_data_toggle),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEFFE;
defparam \WideOr0~0 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_mm_interconnect_0_rsp_demux_009_2 (
	rp_valid,
	always10,
	mem_66_0,
	mem_48_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	rp_valid;
input 	always10;
input 	mem_66_0;
input 	mem_48_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(rp_valid),
	.datab(always10),
	.datac(mem_66_0),
	.datad(mem_48_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hEFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src1_valid~0 (
	.dataa(rp_valid),
	.datab(always10),
	.datac(mem_66_0),
	.datad(mem_48_0),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFFFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_mm_interconnect_0_rsp_mux (
	readdata_0,
	readdata_01,
	readdata_1,
	readdata_11,
	readdata_23,
	readdata_231,
	readdata_22,
	readdata_221,
	readdata_21,
	readdata_211,
	readdata_20,
	readdata_201,
	readdata_19,
	readdata_191,
	readdata_18,
	readdata_181,
	readdata_17,
	readdata_171,
	readdata_16,
	readdata_161,
	read_latency_shift_reg_0,
	mem_84_0,
	mem_66_0,
	read_latency_shift_reg_01,
	out_data_toggle_flopped,
	out_data_toggle_flopped1,
	dreg_0,
	dreg_01,
	out_data_toggle_flopped2,
	dreg_02,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	read_latency_shift_reg_04,
	read_latency_shift_reg_05,
	read_latency_shift_reg_06,
	read_latency_shift_reg_07,
	read_latency_shift_reg_08,
	read_latency_shift_reg_09,
	mem_54_0,
	src0_valid,
	WideOr11,
	av_readdata_pre_0,
	out_payload_0,
	source_addr_1,
	F_iw_0,
	av_readdata_pre_1,
	data_reg_1,
	out_payload_1,
	src_data_1,
	av_readdata_pre_2,
	out_payload_2,
	F_iw_2,
	av_readdata_pre_3,
	data_reg_3,
	out_payload_3,
	src_data_3,
	av_readdata_pre_4,
	data_reg_4,
	out_payload_4,
	src_data_4,
	av_readdata_pre_11,
	data_reg_11,
	out_payload_11,
	src_data_11,
	av_readdata_pre_13,
	data_reg_13,
	out_payload_13,
	src_data_13,
	av_readdata_pre_16,
	av_readdata_pre_12,
	F_iw_12,
	av_readdata_pre_5,
	data_reg_5,
	out_payload_5,
	src_data_5,
	av_readdata_pre_14,
	F_iw_14,
	av_readdata_pre_15,
	data_reg_15,
	out_payload_15,
	src_data_15,
	av_readdata_pre_10,
	F_iw_10,
	av_readdata_pre_9,
	F_iw_9,
	av_readdata_pre_8,
	F_iw_8,
	av_readdata_pre_7,
	out_payload_7,
	F_iw_7,
	av_readdata_pre_6,
	out_payload_6,
	F_iw_6,
	av_readdata_pre_21,
	av_readdata_pre_23,
	av_readdata_pre_22,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	readdata_02,
	av_readdata_pre_01,
	readdata_03,
	readdata_04,
	readdata_05,
	out_valid,
	out_valid1,
	out_data_buffer_0,
	out_data_buffer_01,
	av_readdata_pre_02,
	out_valid2,
	out_data_buffer_02,
	src_data_0,
	readdata_12,
	av_readdata_pre_110,
	readdata_13,
	readdata_14,
	readdata_15,
	out_data_buffer_1,
	out_data_buffer_11,
	av_readdata_pre_111,
	out_data_buffer_12,
	src_data_12,
	src_data_2,
	readdata_2,
	av_readdata_pre_24,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_27,
	out_data_buffer_2,
	av_readdata_pre_25,
	out_data_buffer_21,
	src_data_21,
	readdata_3,
	av_readdata_pre_31,
	readdata_31,
	readdata_32,
	readdata_33,
	readdata_34,
	out_data_buffer_3,
	av_readdata_pre_32,
	out_data_buffer_31,
	src_data_31,
	readdata_4,
	av_readdata_pre_41,
	readdata_41,
	readdata_42,
	readdata_43,
	av_readdata_pre_30,
	out_data_buffer_4,
	av_readdata_pre_42,
	out_data_buffer_41,
	src_data_41,
	readdata_5,
	av_readdata_pre_51,
	src0_valid1,
	readdata_51,
	readdata_52,
	out_data_buffer_5,
	readdata_53,
	av_readdata_pre_52,
	out_data_buffer_51,
	src_data_51,
	readdata_6,
	av_readdata_pre_61,
	readdata_61,
	readdata_62,
	out_data_buffer_6,
	readdata_63,
	av_readdata_pre_62,
	out_data_buffer_61,
	src_data_6,
	readdata_7,
	av_readdata_pre_71,
	readdata_71,
	readdata_72,
	out_data_buffer_7,
	readdata_73,
	av_readdata_pre_72,
	out_data_buffer_71,
	src_data_7,
	src_payload,
	readdata_232,
	out_data_buffer_23,
	src_payload1,
	readdata_222,
	out_data_buffer_22,
	out_data_buffer_221,
	src_payload2,
	readdata_212,
	out_data_buffer_211,
	out_data_buffer_212,
	src_payload3,
	readdata_202,
	out_data_buffer_20,
	out_data_buffer_201,
	src_payload4,
	readdata_192,
	out_data_buffer_19,
	out_data_buffer_191,
	src_payload5,
	readdata_182,
	out_data_buffer_18,
	out_data_buffer_181,
	src_payload6,
	readdata_172,
	out_data_buffer_17,
	out_data_buffer_171,
	src_payload7,
	readdata_162,
	out_data_buffer_16,
	out_data_buffer_161,
	src_payload8,
	readdata_151,
	av_readdata_pre_151,
	readdata_152,
	readdata_153,
	out_data_buffer_15,
	out_data_buffer_151,
	av_readdata_pre_152,
	src_data_151,
	out_data_buffer_14,
	readdata_141,
	av_readdata_pre_141,
	out_data_buffer_141,
	src_data_14,
	av_readdata_pre_131,
	readdata_131,
	out_data_buffer_13,
	out_data_buffer_131,
	src_data_131,
	out_data_buffer_121,
	readdata_121,
	av_readdata_pre_121,
	out_data_buffer_122,
	src_data_121,
	readdata_111,
	av_readdata_pre_112,
	av_readdata_pre_113,
	out_data_buffer_111,
	src_data_111,
	av_readdata_pre_101,
	readdata_10,
	av_readdata_pre_102,
	out_data_buffer_10,
	out_data_buffer_101,
	src_data_10,
	readdata_9,
	av_readdata_pre_91,
	readdata_91,
	readdata_92,
	out_data_buffer_9,
	out_data_buffer_91,
	av_readdata_pre_92,
	src_data_9,
	readdata_8,
	av_readdata_pre_81,
	readdata_81,
	readdata_82,
	out_data_buffer_8,
	av_readdata_pre_82,
	out_data_buffer_81,
	src_data_8)/* synthesis synthesis_greybox=1 */;
input 	readdata_0;
input 	readdata_01;
input 	readdata_1;
input 	readdata_11;
input 	readdata_23;
input 	readdata_231;
input 	readdata_22;
input 	readdata_221;
input 	readdata_21;
input 	readdata_211;
input 	readdata_20;
input 	readdata_201;
input 	readdata_19;
input 	readdata_191;
input 	readdata_18;
input 	readdata_181;
input 	readdata_17;
input 	readdata_171;
input 	readdata_16;
input 	readdata_161;
input 	read_latency_shift_reg_0;
input 	mem_84_0;
input 	mem_66_0;
input 	read_latency_shift_reg_01;
input 	out_data_toggle_flopped;
input 	out_data_toggle_flopped1;
input 	dreg_0;
input 	dreg_01;
input 	out_data_toggle_flopped2;
input 	dreg_02;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	read_latency_shift_reg_04;
input 	read_latency_shift_reg_05;
input 	read_latency_shift_reg_06;
input 	read_latency_shift_reg_07;
input 	read_latency_shift_reg_08;
input 	read_latency_shift_reg_09;
input 	mem_54_0;
input 	src0_valid;
output 	WideOr11;
input 	av_readdata_pre_0;
input 	out_payload_0;
input 	source_addr_1;
input 	F_iw_0;
input 	av_readdata_pre_1;
input 	data_reg_1;
input 	out_payload_1;
output 	src_data_1;
input 	av_readdata_pre_2;
input 	out_payload_2;
input 	F_iw_2;
input 	av_readdata_pre_3;
input 	data_reg_3;
input 	out_payload_3;
output 	src_data_3;
input 	av_readdata_pre_4;
input 	data_reg_4;
input 	out_payload_4;
output 	src_data_4;
input 	av_readdata_pre_11;
input 	data_reg_11;
input 	out_payload_11;
output 	src_data_11;
input 	av_readdata_pre_13;
input 	data_reg_13;
input 	out_payload_13;
output 	src_data_13;
input 	av_readdata_pre_16;
input 	av_readdata_pre_12;
input 	F_iw_12;
input 	av_readdata_pre_5;
input 	data_reg_5;
input 	out_payload_5;
output 	src_data_5;
input 	av_readdata_pre_14;
input 	F_iw_14;
input 	av_readdata_pre_15;
input 	data_reg_15;
input 	out_payload_15;
output 	src_data_15;
input 	av_readdata_pre_10;
input 	F_iw_10;
input 	av_readdata_pre_9;
input 	F_iw_9;
input 	av_readdata_pre_8;
input 	F_iw_8;
input 	av_readdata_pre_7;
input 	out_payload_7;
input 	F_iw_7;
input 	av_readdata_pre_6;
input 	out_payload_6;
input 	F_iw_6;
input 	av_readdata_pre_21;
input 	av_readdata_pre_23;
input 	av_readdata_pre_22;
input 	av_readdata_pre_20;
input 	av_readdata_pre_19;
input 	av_readdata_pre_18;
input 	av_readdata_pre_17;
input 	readdata_02;
input 	av_readdata_pre_01;
input 	readdata_03;
input 	readdata_04;
input 	readdata_05;
input 	out_valid;
input 	out_valid1;
input 	out_data_buffer_0;
input 	out_data_buffer_01;
input 	av_readdata_pre_02;
input 	out_valid2;
input 	out_data_buffer_02;
output 	src_data_0;
input 	readdata_12;
input 	av_readdata_pre_110;
input 	readdata_13;
input 	readdata_14;
input 	readdata_15;
input 	out_data_buffer_1;
input 	out_data_buffer_11;
input 	av_readdata_pre_111;
input 	out_data_buffer_12;
output 	src_data_12;
output 	src_data_2;
input 	readdata_2;
input 	av_readdata_pre_24;
input 	readdata_24;
input 	readdata_25;
input 	readdata_26;
input 	readdata_27;
input 	out_data_buffer_2;
input 	av_readdata_pre_25;
input 	out_data_buffer_21;
output 	src_data_21;
input 	readdata_3;
input 	av_readdata_pre_31;
input 	readdata_31;
input 	readdata_32;
input 	readdata_33;
input 	readdata_34;
input 	out_data_buffer_3;
input 	av_readdata_pre_32;
input 	out_data_buffer_31;
output 	src_data_31;
input 	readdata_4;
input 	av_readdata_pre_41;
input 	readdata_41;
input 	readdata_42;
input 	readdata_43;
input 	av_readdata_pre_30;
input 	out_data_buffer_4;
input 	av_readdata_pre_42;
input 	out_data_buffer_41;
output 	src_data_41;
input 	readdata_5;
input 	av_readdata_pre_51;
input 	src0_valid1;
input 	readdata_51;
input 	readdata_52;
input 	out_data_buffer_5;
input 	readdata_53;
input 	av_readdata_pre_52;
input 	out_data_buffer_51;
output 	src_data_51;
input 	readdata_6;
input 	av_readdata_pre_61;
input 	readdata_61;
input 	readdata_62;
input 	out_data_buffer_6;
input 	readdata_63;
input 	av_readdata_pre_62;
input 	out_data_buffer_61;
output 	src_data_6;
input 	readdata_7;
input 	av_readdata_pre_71;
input 	readdata_71;
input 	readdata_72;
input 	out_data_buffer_7;
input 	readdata_73;
input 	av_readdata_pre_72;
input 	out_data_buffer_71;
output 	src_data_7;
output 	src_payload;
input 	readdata_232;
input 	out_data_buffer_23;
output 	src_payload1;
input 	readdata_222;
input 	out_data_buffer_22;
input 	out_data_buffer_221;
output 	src_payload2;
input 	readdata_212;
input 	out_data_buffer_211;
input 	out_data_buffer_212;
output 	src_payload3;
input 	readdata_202;
input 	out_data_buffer_20;
input 	out_data_buffer_201;
output 	src_payload4;
input 	readdata_192;
input 	out_data_buffer_19;
input 	out_data_buffer_191;
output 	src_payload5;
input 	readdata_182;
input 	out_data_buffer_18;
input 	out_data_buffer_181;
output 	src_payload6;
input 	readdata_172;
input 	out_data_buffer_17;
input 	out_data_buffer_171;
output 	src_payload7;
input 	readdata_162;
input 	out_data_buffer_16;
input 	out_data_buffer_161;
output 	src_payload8;
input 	readdata_151;
input 	av_readdata_pre_151;
input 	readdata_152;
input 	readdata_153;
input 	out_data_buffer_15;
input 	out_data_buffer_151;
input 	av_readdata_pre_152;
output 	src_data_151;
input 	out_data_buffer_14;
input 	readdata_141;
input 	av_readdata_pre_141;
input 	out_data_buffer_141;
output 	src_data_14;
input 	av_readdata_pre_131;
input 	readdata_131;
input 	out_data_buffer_13;
input 	out_data_buffer_131;
output 	src_data_131;
input 	out_data_buffer_121;
input 	readdata_121;
input 	av_readdata_pre_121;
input 	out_data_buffer_122;
output 	src_data_121;
input 	readdata_111;
input 	av_readdata_pre_112;
input 	av_readdata_pre_113;
input 	out_data_buffer_111;
output 	src_data_111;
input 	av_readdata_pre_101;
input 	readdata_10;
input 	av_readdata_pre_102;
input 	out_data_buffer_10;
input 	out_data_buffer_101;
output 	src_data_10;
input 	readdata_9;
input 	av_readdata_pre_91;
input 	readdata_91;
input 	readdata_92;
input 	out_data_buffer_9;
input 	out_data_buffer_91;
input 	av_readdata_pre_92;
output 	src_data_9;
input 	readdata_8;
input 	av_readdata_pre_81;
input 	readdata_81;
input 	readdata_82;
input 	out_data_buffer_8;
input 	av_readdata_pre_82;
input 	out_data_buffer_81;
output 	src_data_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr1~0_combout ;
wire \WideOr1~1_combout ;
wire \WideOr1~2_combout ;
wire \WideOr1~3_combout ;
wire \WideOr1~4_combout ;
wire \src_payload~0_combout ;
wire \src_data[0]~23_combout ;
wire \src_data[0]~24_combout ;
wire \src_data[0]~25_combout ;
wire \src_data[0]~26_combout ;
wire \src_data[0]~27_combout ;
wire \src_data[0]~28_combout ;
wire \src_data[0]~29_combout ;
wire \src_payload~1_combout ;
wire \src_data[1]~31_combout ;
wire \src_data[1]~32_combout ;
wire \src_data[1]~33_combout ;
wire \src_data[1]~34_combout ;
wire \src_data[1]~35_combout ;
wire \src_data[1]~36_combout ;
wire \src_data[1]~37_combout ;
wire \src_payload~2_combout ;
wire \src_data[2]~40_combout ;
wire \src_data[2]~41_combout ;
wire \src_data[2]~42_combout ;
wire \src_data[2]~43_combout ;
wire \src_data[2]~44_combout ;
wire \src_payload~3_combout ;
wire \src_data[3]~46_combout ;
wire \src_data[3]~47_combout ;
wire \src_data[3]~48_combout ;
wire \src_data[3]~49_combout ;
wire \src_data[3]~50_combout ;
wire \src_data[3]~51_combout ;
wire \src_payload~4_combout ;
wire \src_data[4]~53_combout ;
wire \src_data[4]~54_combout ;
wire \src_data[4]~55_combout ;
wire \src_data[4]~56_combout ;
wire \src_data[4]~57_combout ;
wire \src_data[4]~114_combout ;
wire \src_data[5]~59_combout ;
wire \src_data[5]~60_combout ;
wire \src_data[5]~61_combout ;
wire \src_data[5]~62_combout ;
wire \src_data[5]~63_combout ;
wire \src_data[5]~115_combout ;
wire \src_data[6]~65_combout ;
wire \src_data[6]~66_combout ;
wire \src_data[6]~67_combout ;
wire \src_data[6]~68_combout ;
wire \src_data[6]~69_combout ;
wire \src_data[6]~116_combout ;
wire \src_data[7]~71_combout ;
wire \src_data[7]~72_combout ;
wire \src_data[7]~73_combout ;
wire \src_data[7]~74_combout ;
wire \src_data[7]~75_combout ;
wire \src_data[7]~117_combout ;
wire \src_payload~6_combout ;
wire \src_payload~7_combout ;
wire \src_payload~8_combout ;
wire \src_payload~10_combout ;
wire \src_payload~11_combout ;
wire \src_payload~12_combout ;
wire \src_payload~13_combout ;
wire \src_payload~15_combout ;
wire \src_payload~16_combout ;
wire \src_payload~17_combout ;
wire \src_payload~18_combout ;
wire \src_payload~20_combout ;
wire \src_payload~21_combout ;
wire \src_payload~22_combout ;
wire \src_payload~23_combout ;
wire \src_payload~25_combout ;
wire \src_payload~26_combout ;
wire \src_payload~27_combout ;
wire \src_payload~28_combout ;
wire \src_payload~30_combout ;
wire \src_payload~31_combout ;
wire \src_payload~32_combout ;
wire \src_payload~33_combout ;
wire \src_payload~35_combout ;
wire \src_payload~36_combout ;
wire \src_payload~37_combout ;
wire \src_payload~38_combout ;
wire \src_payload~40_combout ;
wire \src_payload~41_combout ;
wire \src_payload~42_combout ;
wire \src_payload~43_combout ;
wire \src_data[15]~77_combout ;
wire \src_data[15]~78_combout ;
wire \src_data[15]~79_combout ;
wire \src_data[15]~80_combout ;
wire \src_data[15]~81_combout ;
wire \src_data[14]~83_combout ;
wire \src_data[14]~84_combout ;
wire \src_data[14]~118_combout ;
wire \src_payload~45_combout ;
wire \src_data[13]~86_combout ;
wire \src_data[13]~87_combout ;
wire \src_data[13]~88_combout ;
wire \src_data[12]~90_combout ;
wire \src_data[12]~91_combout ;
wire \src_data[12]~119_combout ;
wire \src_data[11]~93_combout ;
wire \src_data[11]~94_combout ;
wire \src_data[11]~95_combout ;
wire \src_data[11]~120_combout ;
wire \src_data[10]~97_combout ;
wire \src_data[10]~98_combout ;
wire \src_data[10]~99_combout ;
wire \src_data[10]~100_combout ;
wire \src_data[9]~102_combout ;
wire \src_data[9]~103_combout ;
wire \src_data[9]~104_combout ;
wire \src_data[9]~105_combout ;
wire \src_data[9]~106_combout ;
wire \src_data[8]~108_combout ;
wire \src_data[8]~109_combout ;
wire \src_data[8]~110_combout ;
wire \src_data[8]~111_combout ;
wire \src_data[8]~112_combout ;
wire \src_data[8]~121_combout ;


cycloneive_lcell_comb WideOr1(
	.dataa(\WideOr1~4_combout ),
	.datab(read_latency_shift_reg_08),
	.datac(read_latency_shift_reg_09),
	.datad(src0_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hBFFF;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~16 (
	.dataa(mem_54_0),
	.datab(data_reg_1),
	.datac(out_payload_1),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(src_data_1),
	.cout());
defparam \src_data[1]~16 .lut_mask = 16'hFEFF;
defparam \src_data[1]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~17 (
	.dataa(mem_54_0),
	.datab(data_reg_3),
	.datac(out_payload_3),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(src_data_3),
	.cout());
defparam \src_data[3]~17 .lut_mask = 16'hFEFF;
defparam \src_data[3]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~18 (
	.dataa(mem_54_0),
	.datab(data_reg_4),
	.datac(out_payload_4),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(src_data_4),
	.cout());
defparam \src_data[4]~18 .lut_mask = 16'hFEFF;
defparam \src_data[4]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~19 (
	.dataa(mem_54_0),
	.datab(data_reg_11),
	.datac(out_payload_11),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(src_data_11),
	.cout());
defparam \src_data[11]~19 .lut_mask = 16'hFEFF;
defparam \src_data[11]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~20 (
	.dataa(mem_54_0),
	.datab(data_reg_13),
	.datac(out_payload_13),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(src_data_13),
	.cout());
defparam \src_data[13]~20 .lut_mask = 16'hFEFF;
defparam \src_data[13]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~21 (
	.dataa(mem_54_0),
	.datab(data_reg_5),
	.datac(out_payload_5),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(src_data_5),
	.cout());
defparam \src_data[5]~21 .lut_mask = 16'hFEFF;
defparam \src_data[5]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~22 (
	.dataa(mem_54_0),
	.datab(data_reg_15),
	.datac(out_payload_15),
	.datad(source_addr_1),
	.cin(gnd),
	.combout(src_data_15),
	.cout());
defparam \src_data[15]~22 .lut_mask = 16'hFEFF;
defparam \src_data[15]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~30 (
	.dataa(\src_data[0]~26_combout ),
	.datab(\src_data[0]~29_combout ),
	.datac(src0_valid),
	.datad(F_iw_0),
	.cin(gnd),
	.combout(src_data_0),
	.cout());
defparam \src_data[0]~30 .lut_mask = 16'hFFFE;
defparam \src_data[0]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~38 (
	.dataa(\src_data[1]~34_combout ),
	.datab(\src_data[1]~37_combout ),
	.datac(src0_valid),
	.datad(src_data_1),
	.cin(gnd),
	.combout(src_data_12),
	.cout());
defparam \src_data[1]~38 .lut_mask = 16'hFFFE;
defparam \src_data[1]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~39 (
	.dataa(src0_valid),
	.datab(F_iw_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_2),
	.cout());
defparam \src_data[2]~39 .lut_mask = 16'hEEEE;
defparam \src_data[2]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~45 (
	.dataa(\src_data[2]~43_combout ),
	.datab(\src_data[2]~44_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_21),
	.cin(gnd),
	.combout(src_data_21),
	.cout());
defparam \src_data[2]~45 .lut_mask = 16'hFFFE;
defparam \src_data[2]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~52 (
	.dataa(\src_data[3]~51_combout ),
	.datab(src0_valid),
	.datac(src_data_3),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_31),
	.cout());
defparam \src_data[3]~52 .lut_mask = 16'hFEFE;
defparam \src_data[3]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~58 (
	.dataa(\src_data[4]~56_combout ),
	.datab(\src_data[4]~114_combout ),
	.datac(src0_valid),
	.datad(src_data_4),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[4]~58 .lut_mask = 16'hFFFE;
defparam \src_data[4]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~64 (
	.dataa(\src_data[5]~62_combout ),
	.datab(\src_data[5]~115_combout ),
	.datac(src0_valid),
	.datad(src_data_5),
	.cin(gnd),
	.combout(src_data_51),
	.cout());
defparam \src_data[5]~64 .lut_mask = 16'hFFFE;
defparam \src_data[5]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~70 (
	.dataa(\src_data[6]~68_combout ),
	.datab(\src_data[6]~116_combout ),
	.datac(src0_valid),
	.datad(F_iw_6),
	.cin(gnd),
	.combout(src_data_6),
	.cout());
defparam \src_data[6]~70 .lut_mask = 16'hFFFE;
defparam \src_data[6]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~76 (
	.dataa(\src_data[7]~74_combout ),
	.datab(\src_data[7]~117_combout ),
	.datac(src0_valid),
	.datad(F_iw_7),
	.cin(gnd),
	.combout(src_data_7),
	.cout());
defparam \src_data[7]~76 .lut_mask = 16'hFFFE;
defparam \src_data[7]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(source_addr_1),
	.datab(src0_valid),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(\src_payload~8_combout ),
	.datab(source_addr_1),
	.datac(src0_valid),
	.datad(out_payload_7),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hFFFE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(\src_payload~10_combout ),
	.datab(\src_payload~13_combout ),
	.datac(out_payload_6),
	.datad(src_payload),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hFFFE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(\src_payload~15_combout ),
	.datab(\src_payload~18_combout ),
	.datac(out_payload_5),
	.datad(src_payload),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hFFFE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~24 (
	.dataa(\src_payload~20_combout ),
	.datab(\src_payload~23_combout ),
	.datac(out_payload_4),
	.datad(src_payload),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hFFFE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~29 (
	.dataa(\src_payload~25_combout ),
	.datab(\src_payload~28_combout ),
	.datac(out_payload_3),
	.datad(src_payload),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hFFFE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~34 (
	.dataa(\src_payload~30_combout ),
	.datab(\src_payload~33_combout ),
	.datac(out_payload_2),
	.datad(src_payload),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~34 .lut_mask = 16'hFFFE;
defparam \src_payload~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~39 (
	.dataa(\src_payload~35_combout ),
	.datab(\src_payload~38_combout ),
	.datac(out_payload_1),
	.datad(src_payload),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~39 .lut_mask = 16'hFFFE;
defparam \src_payload~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~44 (
	.dataa(\src_payload~40_combout ),
	.datab(\src_payload~43_combout ),
	.datac(out_payload_0),
	.datad(src_payload),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~44 .lut_mask = 16'hFFFE;
defparam \src_payload~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~82 (
	.dataa(\src_data[15]~80_combout ),
	.datab(\src_data[15]~81_combout ),
	.datac(src0_valid),
	.datad(src_data_15),
	.cin(gnd),
	.combout(src_data_151),
	.cout());
defparam \src_data[15]~82 .lut_mask = 16'hFFFE;
defparam \src_data[15]~82 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~85 (
	.dataa(\src_data[14]~83_combout ),
	.datab(\src_data[14]~118_combout ),
	.datac(src0_valid),
	.datad(F_iw_14),
	.cin(gnd),
	.combout(src_data_14),
	.cout());
defparam \src_data[14]~85 .lut_mask = 16'hFFFE;
defparam \src_data[14]~85 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~89 (
	.dataa(\src_payload~45_combout ),
	.datab(\src_data[13]~88_combout ),
	.datac(src0_valid),
	.datad(src_data_13),
	.cin(gnd),
	.combout(src_data_131),
	.cout());
defparam \src_data[13]~89 .lut_mask = 16'hFFFE;
defparam \src_data[13]~89 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~92 (
	.dataa(\src_data[12]~90_combout ),
	.datab(\src_data[12]~119_combout ),
	.datac(src0_valid),
	.datad(F_iw_12),
	.cin(gnd),
	.combout(src_data_121),
	.cout());
defparam \src_data[12]~92 .lut_mask = 16'hFFFE;
defparam \src_data[12]~92 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~96 (
	.dataa(\src_data[11]~94_combout ),
	.datab(\src_data[11]~120_combout ),
	.datac(src0_valid),
	.datad(src_data_11),
	.cin(gnd),
	.combout(src_data_111),
	.cout());
defparam \src_data[11]~96 .lut_mask = 16'hFFFE;
defparam \src_data[11]~96 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~101 (
	.dataa(\src_data[10]~97_combout ),
	.datab(\src_data[10]~100_combout ),
	.datac(src0_valid),
	.datad(F_iw_10),
	.cin(gnd),
	.combout(src_data_10),
	.cout());
defparam \src_data[10]~101 .lut_mask = 16'hFFFE;
defparam \src_data[10]~101 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~107 (
	.dataa(\src_data[9]~105_combout ),
	.datab(\src_data[9]~106_combout ),
	.datac(src0_valid),
	.datad(F_iw_9),
	.cin(gnd),
	.combout(src_data_9),
	.cout());
defparam \src_data[9]~107 .lut_mask = 16'hFFFE;
defparam \src_data[9]~107 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~113 (
	.dataa(\src_data[8]~111_combout ),
	.datab(\src_data[8]~121_combout ),
	.datac(src0_valid),
	.datad(F_iw_8),
	.cin(gnd),
	.combout(src_data_8),
	.cout());
defparam \src_data[8]~113 .lut_mask = 16'hFFFE;
defparam \src_data[8]~113 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~0 (
	.dataa(mem_84_0),
	.datab(mem_66_0),
	.datac(read_latency_shift_reg_01),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hEFFF;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~1 (
	.dataa(out_data_toggle_flopped),
	.datab(out_data_toggle_flopped1),
	.datac(dreg_0),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\WideOr1~1_combout ),
	.cout());
defparam \WideOr1~1 .lut_mask = 16'h6996;
defparam \WideOr1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~2 (
	.dataa(out_data_toggle_flopped2),
	.datab(dreg_02),
	.datac(read_latency_shift_reg_02),
	.datad(read_latency_shift_reg_03),
	.cin(gnd),
	.combout(\WideOr1~2_combout ),
	.cout());
defparam \WideOr1~2 .lut_mask = 16'h6FFF;
defparam \WideOr1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~3 (
	.dataa(read_latency_shift_reg_04),
	.datab(read_latency_shift_reg_05),
	.datac(read_latency_shift_reg_06),
	.datad(read_latency_shift_reg_07),
	.cin(gnd),
	.combout(\WideOr1~3_combout ),
	.cout());
defparam \WideOr1~3 .lut_mask = 16'h7FFF;
defparam \WideOr1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~4 (
	.dataa(\WideOr1~0_combout ),
	.datab(\WideOr1~1_combout ),
	.datac(\WideOr1~2_combout ),
	.datad(\WideOr1~3_combout ),
	.cin(gnd),
	.combout(\WideOr1~4_combout ),
	.cout());
defparam \WideOr1~4 .lut_mask = 16'hFFFE;
defparam \WideOr1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_0),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\src_payload~0_combout ),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEFFF;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~23 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_02),
	.datac(readdata_02),
	.datad(av_readdata_pre_01),
	.cin(gnd),
	.combout(\src_data[0]~23_combout ),
	.cout());
defparam \src_data[0]~23 .lut_mask = 16'hFFFE;
defparam \src_data[0]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~24 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(readdata_03),
	.datad(readdata_04),
	.cin(gnd),
	.combout(\src_data[0]~24_combout ),
	.cout());
defparam \src_data[0]~24 .lut_mask = 16'hFFFE;
defparam \src_data[0]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~25 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_0),
	.datad(readdata_05),
	.cin(gnd),
	.combout(\src_data[0]~25_combout ),
	.cout());
defparam \src_data[0]~25 .lut_mask = 16'hFFFE;
defparam \src_data[0]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~26 (
	.dataa(\src_payload~0_combout ),
	.datab(\src_data[0]~23_combout ),
	.datac(\src_data[0]~24_combout ),
	.datad(\src_data[0]~25_combout ),
	.cin(gnd),
	.combout(\src_data[0]~26_combout ),
	.cout());
defparam \src_data[0]~26 .lut_mask = 16'hFFFE;
defparam \src_data[0]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~27 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_0),
	.datad(out_data_buffer_01),
	.cin(gnd),
	.combout(\src_data[0]~27_combout ),
	.cout());
defparam \src_data[0]~27 .lut_mask = 16'hFFFE;
defparam \src_data[0]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~28 (
	.dataa(read_latency_shift_reg_09),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_01),
	.datad(av_readdata_pre_02),
	.cin(gnd),
	.combout(\src_data[0]~28_combout ),
	.cout());
defparam \src_data[0]~28 .lut_mask = 16'hFFFE;
defparam \src_data[0]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~29 (
	.dataa(\src_data[0]~27_combout ),
	.datab(\src_data[0]~28_combout ),
	.datac(out_valid2),
	.datad(out_data_buffer_02),
	.cin(gnd),
	.combout(\src_data[0]~29_combout ),
	.cout());
defparam \src_data[0]~29 .lut_mask = 16'hFFFE;
defparam \src_data[0]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_1),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\src_payload~1_combout ),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEFFF;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~31 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_02),
	.datac(readdata_12),
	.datad(av_readdata_pre_110),
	.cin(gnd),
	.combout(\src_data[1]~31_combout ),
	.cout());
defparam \src_data[1]~31 .lut_mask = 16'hFFFE;
defparam \src_data[1]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~32 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(readdata_13),
	.datad(readdata_14),
	.cin(gnd),
	.combout(\src_data[1]~32_combout ),
	.cout());
defparam \src_data[1]~32 .lut_mask = 16'hFFFE;
defparam \src_data[1]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~33 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_1),
	.datad(readdata_15),
	.cin(gnd),
	.combout(\src_data[1]~33_combout ),
	.cout());
defparam \src_data[1]~33 .lut_mask = 16'hFFFE;
defparam \src_data[1]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~34 (
	.dataa(\src_payload~1_combout ),
	.datab(\src_data[1]~31_combout ),
	.datac(\src_data[1]~32_combout ),
	.datad(\src_data[1]~33_combout ),
	.cin(gnd),
	.combout(\src_data[1]~34_combout ),
	.cout());
defparam \src_data[1]~34 .lut_mask = 16'hFFFE;
defparam \src_data[1]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~35 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_1),
	.datad(out_data_buffer_11),
	.cin(gnd),
	.combout(\src_data[1]~35_combout ),
	.cout());
defparam \src_data[1]~35 .lut_mask = 16'hFFFE;
defparam \src_data[1]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~36 (
	.dataa(read_latency_shift_reg_09),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_11),
	.datad(av_readdata_pre_111),
	.cin(gnd),
	.combout(\src_data[1]~36_combout ),
	.cout());
defparam \src_data[1]~36 .lut_mask = 16'hFFFE;
defparam \src_data[1]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~37 (
	.dataa(\src_data[1]~35_combout ),
	.datab(\src_data[1]~36_combout ),
	.datac(out_valid2),
	.datad(out_data_buffer_12),
	.cin(gnd),
	.combout(\src_data[1]~37_combout ),
	.cout());
defparam \src_data[1]~37 .lut_mask = 16'hFFFE;
defparam \src_data[1]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_2),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\src_payload~2_combout ),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEFFF;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~40 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_02),
	.datac(readdata_2),
	.datad(av_readdata_pre_24),
	.cin(gnd),
	.combout(\src_data[2]~40_combout ),
	.cout());
defparam \src_data[2]~40 .lut_mask = 16'hFFFE;
defparam \src_data[2]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~41 (
	.dataa(read_latency_shift_reg_04),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_24),
	.datad(readdata_25),
	.cin(gnd),
	.combout(\src_data[2]~41_combout ),
	.cout());
defparam \src_data[2]~41 .lut_mask = 16'hFFFE;
defparam \src_data[2]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~42 (
	.dataa(read_latency_shift_reg_06),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_26),
	.datad(readdata_27),
	.cin(gnd),
	.combout(\src_data[2]~42_combout ),
	.cout());
defparam \src_data[2]~42 .lut_mask = 16'hFFFE;
defparam \src_data[2]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~43 (
	.dataa(\src_payload~2_combout ),
	.datab(\src_data[2]~40_combout ),
	.datac(\src_data[2]~41_combout ),
	.datad(\src_data[2]~42_combout ),
	.cin(gnd),
	.combout(\src_data[2]~43_combout ),
	.cout());
defparam \src_data[2]~43 .lut_mask = 16'hFFFE;
defparam \src_data[2]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~44 (
	.dataa(read_latency_shift_reg_09),
	.datab(out_valid1),
	.datac(out_data_buffer_2),
	.datad(av_readdata_pre_25),
	.cin(gnd),
	.combout(\src_data[2]~44_combout ),
	.cout());
defparam \src_data[2]~44 .lut_mask = 16'hFFFE;
defparam \src_data[2]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_3),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\src_payload~3_combout ),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEFFF;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~46 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_02),
	.datac(readdata_3),
	.datad(av_readdata_pre_31),
	.cin(gnd),
	.combout(\src_data[3]~46_combout ),
	.cout());
defparam \src_data[3]~46 .lut_mask = 16'hFFFE;
defparam \src_data[3]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~47 (
	.dataa(read_latency_shift_reg_04),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_31),
	.datad(readdata_32),
	.cin(gnd),
	.combout(\src_data[3]~47_combout ),
	.cout());
defparam \src_data[3]~47 .lut_mask = 16'hFFFE;
defparam \src_data[3]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~48 (
	.dataa(read_latency_shift_reg_06),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_33),
	.datad(readdata_34),
	.cin(gnd),
	.combout(\src_data[3]~48_combout ),
	.cout());
defparam \src_data[3]~48 .lut_mask = 16'hFFFE;
defparam \src_data[3]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~49 (
	.dataa(\src_payload~3_combout ),
	.datab(\src_data[3]~46_combout ),
	.datac(\src_data[3]~47_combout ),
	.datad(\src_data[3]~48_combout ),
	.cin(gnd),
	.combout(\src_data[3]~49_combout ),
	.cout());
defparam \src_data[3]~49 .lut_mask = 16'hFFFE;
defparam \src_data[3]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~50 (
	.dataa(read_latency_shift_reg_09),
	.datab(out_valid1),
	.datac(out_data_buffer_3),
	.datad(av_readdata_pre_32),
	.cin(gnd),
	.combout(\src_data[3]~50_combout ),
	.cout());
defparam \src_data[3]~50 .lut_mask = 16'hFFFE;
defparam \src_data[3]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~51 (
	.dataa(\src_data[3]~49_combout ),
	.datab(\src_data[3]~50_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_31),
	.cin(gnd),
	.combout(\src_data[3]~51_combout ),
	.cout());
defparam \src_data[3]~51 .lut_mask = 16'hFFFE;
defparam \src_data[3]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_4),
	.datac(mem_84_0),
	.datad(mem_66_0),
	.cin(gnd),
	.combout(\src_payload~4_combout ),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEFFF;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~53 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_02),
	.datac(readdata_4),
	.datad(av_readdata_pre_41),
	.cin(gnd),
	.combout(\src_data[4]~53_combout ),
	.cout());
defparam \src_data[4]~53 .lut_mask = 16'hFFFE;
defparam \src_data[4]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~54 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_41),
	.datad(readdata_42),
	.cin(gnd),
	.combout(\src_data[4]~54_combout ),
	.cout());
defparam \src_data[4]~54 .lut_mask = 16'hFFFE;
defparam \src_data[4]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~55 (
	.dataa(read_latency_shift_reg_08),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_43),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\src_data[4]~55_combout ),
	.cout());
defparam \src_data[4]~55 .lut_mask = 16'hFFFE;
defparam \src_data[4]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~56 (
	.dataa(\src_payload~4_combout ),
	.datab(\src_data[4]~53_combout ),
	.datac(\src_data[4]~54_combout ),
	.datad(\src_data[4]~55_combout ),
	.cin(gnd),
	.combout(\src_data[4]~56_combout ),
	.cout());
defparam \src_data[4]~56 .lut_mask = 16'hFFFE;
defparam \src_data[4]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~57 (
	.dataa(read_latency_shift_reg_09),
	.datab(out_valid1),
	.datac(out_data_buffer_4),
	.datad(av_readdata_pre_42),
	.cin(gnd),
	.combout(\src_data[4]~57_combout ),
	.cout());
defparam \src_data[4]~57 .lut_mask = 16'hFFFE;
defparam \src_data[4]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~114 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_01),
	.datac(\src_data[4]~57_combout ),
	.datad(out_data_buffer_41),
	.cin(gnd),
	.combout(\src_data[4]~114_combout ),
	.cout());
defparam \src_data[4]~114 .lut_mask = 16'hFFF6;
defparam \src_data[4]~114 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~59 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_02),
	.datac(readdata_5),
	.datad(av_readdata_pre_51),
	.cin(gnd),
	.combout(\src_data[5]~59_combout ),
	.cout());
defparam \src_data[5]~59 .lut_mask = 16'hFFFE;
defparam \src_data[5]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~60 (
	.dataa(\src_data[5]~59_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[5]~60_combout ),
	.cout());
defparam \src_data[5]~60 .lut_mask = 16'hFEFE;
defparam \src_data[5]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~61 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_51),
	.datad(readdata_52),
	.cin(gnd),
	.combout(\src_data[5]~61_combout ),
	.cout());
defparam \src_data[5]~61 .lut_mask = 16'hFFFE;
defparam \src_data[5]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~62 (
	.dataa(\src_data[5]~60_combout ),
	.datab(\src_data[5]~61_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_5),
	.cin(gnd),
	.combout(\src_data[5]~62_combout ),
	.cout());
defparam \src_data[5]~62 .lut_mask = 16'hFFFE;
defparam \src_data[5]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~63 (
	.dataa(read_latency_shift_reg_09),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_53),
	.datad(av_readdata_pre_52),
	.cin(gnd),
	.combout(\src_data[5]~63_combout ),
	.cout());
defparam \src_data[5]~63 .lut_mask = 16'hFFFE;
defparam \src_data[5]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~115 (
	.dataa(out_data_toggle_flopped1),
	.datab(dreg_0),
	.datac(\src_data[5]~63_combout ),
	.datad(out_data_buffer_51),
	.cin(gnd),
	.combout(\src_data[5]~115_combout ),
	.cout());
defparam \src_data[5]~115 .lut_mask = 16'hFFF6;
defparam \src_data[5]~115 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~65 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_02),
	.datac(readdata_6),
	.datad(av_readdata_pre_61),
	.cin(gnd),
	.combout(\src_data[6]~65_combout ),
	.cout());
defparam \src_data[6]~65 .lut_mask = 16'hFFFE;
defparam \src_data[6]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~66 (
	.dataa(\src_data[6]~65_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[6]~66_combout ),
	.cout());
defparam \src_data[6]~66 .lut_mask = 16'hFEFE;
defparam \src_data[6]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~67 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_61),
	.datad(readdata_62),
	.cin(gnd),
	.combout(\src_data[6]~67_combout ),
	.cout());
defparam \src_data[6]~67 .lut_mask = 16'hFFFE;
defparam \src_data[6]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~68 (
	.dataa(\src_data[6]~66_combout ),
	.datab(\src_data[6]~67_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_6),
	.cin(gnd),
	.combout(\src_data[6]~68_combout ),
	.cout());
defparam \src_data[6]~68 .lut_mask = 16'hFFFE;
defparam \src_data[6]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~69 (
	.dataa(read_latency_shift_reg_09),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_63),
	.datad(av_readdata_pre_62),
	.cin(gnd),
	.combout(\src_data[6]~69_combout ),
	.cout());
defparam \src_data[6]~69 .lut_mask = 16'hFFFE;
defparam \src_data[6]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~116 (
	.dataa(out_data_toggle_flopped1),
	.datab(dreg_0),
	.datac(\src_data[6]~69_combout ),
	.datad(out_data_buffer_61),
	.cin(gnd),
	.combout(\src_data[6]~116_combout ),
	.cout());
defparam \src_data[6]~116 .lut_mask = 16'hFFF6;
defparam \src_data[6]~116 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~71 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_02),
	.datac(readdata_7),
	.datad(av_readdata_pre_71),
	.cin(gnd),
	.combout(\src_data[7]~71_combout ),
	.cout());
defparam \src_data[7]~71 .lut_mask = 16'hFFFE;
defparam \src_data[7]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~72 (
	.dataa(\src_data[7]~71_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[7]~72_combout ),
	.cout());
defparam \src_data[7]~72 .lut_mask = 16'hFEFE;
defparam \src_data[7]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~73 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_71),
	.datad(readdata_72),
	.cin(gnd),
	.combout(\src_data[7]~73_combout ),
	.cout());
defparam \src_data[7]~73 .lut_mask = 16'hFFFE;
defparam \src_data[7]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~74 (
	.dataa(\src_data[7]~72_combout ),
	.datab(\src_data[7]~73_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_7),
	.cin(gnd),
	.combout(\src_data[7]~74_combout ),
	.cout());
defparam \src_data[7]~74 .lut_mask = 16'hFFFE;
defparam \src_data[7]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~75 (
	.dataa(read_latency_shift_reg_09),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_73),
	.datad(av_readdata_pre_72),
	.cin(gnd),
	.combout(\src_data[7]~75_combout ),
	.cout());
defparam \src_data[7]~75 .lut_mask = 16'hFFFE;
defparam \src_data[7]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~117 (
	.dataa(out_data_toggle_flopped1),
	.datab(dreg_0),
	.datac(\src_data[7]~75_combout ),
	.datad(out_data_buffer_71),
	.cin(gnd),
	.combout(\src_data[7]~117_combout ),
	.cout());
defparam \src_data[7]~117 .lut_mask = 16'hFFF6;
defparam \src_data[7]~117 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_23),
	.datad(readdata_232),
	.cin(gnd),
	.combout(\src_payload~6_combout ),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hFFFE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(out_valid1),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_231),
	.datad(out_data_buffer_23),
	.cin(gnd),
	.combout(\src_payload~7_combout ),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hFFFE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(\src_payload~6_combout ),
	.datab(\src_payload~7_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_23),
	.cin(gnd),
	.combout(\src_payload~8_combout ),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hFFFE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(read_latency_shift_reg_07),
	.datab(readdata_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~10_combout ),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_221),
	.datad(readdata_222),
	.cin(gnd),
	.combout(\src_payload~11_combout ),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hFFFE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_22),
	.datad(out_data_buffer_221),
	.cin(gnd),
	.combout(\src_payload~12_combout ),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hFFFE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(\src_payload~11_combout ),
	.datab(\src_payload~12_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_22),
	.cin(gnd),
	.combout(\src_payload~13_combout ),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hFFFE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(read_latency_shift_reg_07),
	.datab(readdata_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~15_combout ),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_211),
	.datad(readdata_212),
	.cin(gnd),
	.combout(\src_payload~16_combout ),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hFFFE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_211),
	.datad(out_data_buffer_212),
	.cin(gnd),
	.combout(\src_payload~17_combout ),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hFFFE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(\src_payload~16_combout ),
	.datab(\src_payload~17_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_21),
	.cin(gnd),
	.combout(\src_payload~18_combout ),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hFFFE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(read_latency_shift_reg_07),
	.datab(readdata_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~20_combout ),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~21 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_201),
	.datad(readdata_202),
	.cin(gnd),
	.combout(\src_payload~21_combout ),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hFFFE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~22 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_20),
	.datad(out_data_buffer_201),
	.cin(gnd),
	.combout(\src_payload~22_combout ),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hFFFE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~23 (
	.dataa(\src_payload~21_combout ),
	.datab(\src_payload~22_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_20),
	.cin(gnd),
	.combout(\src_payload~23_combout ),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hFFFE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~25 (
	.dataa(read_latency_shift_reg_08),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_19),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\src_payload~25_combout ),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hFFFE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~26 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_191),
	.datad(readdata_192),
	.cin(gnd),
	.combout(\src_payload~26_combout ),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hFFFE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~27 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_19),
	.datad(out_data_buffer_191),
	.cin(gnd),
	.combout(\src_payload~27_combout ),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hFFFE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~28 (
	.dataa(\src_payload~26_combout ),
	.datab(\src_payload~27_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_19),
	.cin(gnd),
	.combout(\src_payload~28_combout ),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hFFFE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~30 (
	.dataa(read_latency_shift_reg_07),
	.datab(readdata_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~30_combout ),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~31 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_181),
	.datad(readdata_182),
	.cin(gnd),
	.combout(\src_payload~31_combout ),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hFFFE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~32 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_18),
	.datad(out_data_buffer_181),
	.cin(gnd),
	.combout(\src_payload~32_combout ),
	.cout());
defparam \src_payload~32 .lut_mask = 16'hFFFE;
defparam \src_payload~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~33 (
	.dataa(\src_payload~31_combout ),
	.datab(\src_payload~32_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_18),
	.cin(gnd),
	.combout(\src_payload~33_combout ),
	.cout());
defparam \src_payload~33 .lut_mask = 16'hFFFE;
defparam \src_payload~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~35 (
	.dataa(read_latency_shift_reg_07),
	.datab(readdata_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~35_combout ),
	.cout());
defparam \src_payload~35 .lut_mask = 16'hEEEE;
defparam \src_payload~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~36 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_171),
	.datad(readdata_172),
	.cin(gnd),
	.combout(\src_payload~36_combout ),
	.cout());
defparam \src_payload~36 .lut_mask = 16'hFFFE;
defparam \src_payload~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~37 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_17),
	.datad(out_data_buffer_171),
	.cin(gnd),
	.combout(\src_payload~37_combout ),
	.cout());
defparam \src_payload~37 .lut_mask = 16'hFFFE;
defparam \src_payload~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~38 (
	.dataa(\src_payload~36_combout ),
	.datab(\src_payload~37_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_17),
	.cin(gnd),
	.combout(\src_payload~38_combout ),
	.cout());
defparam \src_payload~38 .lut_mask = 16'hFFFE;
defparam \src_payload~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~40 (
	.dataa(read_latency_shift_reg_08),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_16),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\src_payload~40_combout ),
	.cout());
defparam \src_payload~40 .lut_mask = 16'hFFFE;
defparam \src_payload~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~41 (
	.dataa(read_latency_shift_reg_05),
	.datab(read_latency_shift_reg_06),
	.datac(readdata_161),
	.datad(readdata_162),
	.cin(gnd),
	.combout(\src_payload~41_combout ),
	.cout());
defparam \src_payload~41 .lut_mask = 16'hFFFE;
defparam \src_payload~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~42 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_16),
	.datad(out_data_buffer_161),
	.cin(gnd),
	.combout(\src_payload~42_combout ),
	.cout());
defparam \src_payload~42 .lut_mask = 16'hFFFE;
defparam \src_payload~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~43 (
	.dataa(\src_payload~41_combout ),
	.datab(\src_payload~42_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_16),
	.cin(gnd),
	.combout(\src_payload~43_combout ),
	.cout());
defparam \src_payload~43 .lut_mask = 16'hFFFE;
defparam \src_payload~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~77 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_151),
	.datad(av_readdata_pre_151),
	.cin(gnd),
	.combout(\src_data[15]~77_combout ),
	.cout());
defparam \src_data[15]~77 .lut_mask = 16'hFFFE;
defparam \src_data[15]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~78 (
	.dataa(\src_data[15]~77_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_15),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[15]~78_combout ),
	.cout());
defparam \src_data[15]~78 .lut_mask = 16'hFEFE;
defparam \src_data[15]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~79 (
	.dataa(read_latency_shift_reg_06),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_152),
	.datad(readdata_153),
	.cin(gnd),
	.combout(\src_data[15]~79_combout ),
	.cout());
defparam \src_data[15]~79 .lut_mask = 16'hFFFE;
defparam \src_data[15]~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~80 (
	.dataa(\src_data[15]~78_combout ),
	.datab(\src_data[15]~79_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_15),
	.cin(gnd),
	.combout(\src_data[15]~80_combout ),
	.cout());
defparam \src_data[15]~80 .lut_mask = 16'hFFFE;
defparam \src_data[15]~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~81 (
	.dataa(read_latency_shift_reg_09),
	.datab(out_valid1),
	.datac(out_data_buffer_151),
	.datad(av_readdata_pre_152),
	.cin(gnd),
	.combout(\src_data[15]~81_combout ),
	.cout());
defparam \src_data[15]~81 .lut_mask = 16'hFFFE;
defparam \src_data[15]~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~83 (
	.dataa(src0_valid1),
	.datab(out_valid),
	.datac(out_data_buffer_14),
	.datad(av_readdata_pre_14),
	.cin(gnd),
	.combout(\src_data[14]~83_combout ),
	.cout());
defparam \src_data[14]~83 .lut_mask = 16'hFFFE;
defparam \src_data[14]~83 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~84 (
	.dataa(read_latency_shift_reg_09),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_141),
	.datad(av_readdata_pre_141),
	.cin(gnd),
	.combout(\src_data[14]~84_combout ),
	.cout());
defparam \src_data[14]~84 .lut_mask = 16'hFFFE;
defparam \src_data[14]~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~118 (
	.dataa(out_data_toggle_flopped1),
	.datab(dreg_0),
	.datac(\src_data[14]~84_combout ),
	.datad(out_data_buffer_141),
	.cin(gnd),
	.combout(\src_data[14]~118_combout ),
	.cout());
defparam \src_data[14]~118 .lut_mask = 16'hFFF6;
defparam \src_data[14]~118 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~45 (
	.dataa(read_latency_shift_reg_09),
	.datab(av_readdata_pre_131),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~45_combout ),
	.cout());
defparam \src_payload~45 .lut_mask = 16'hEEEE;
defparam \src_payload~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~86 (
	.dataa(read_latency_shift_reg_08),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_131),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\src_data[13]~86_combout ),
	.cout());
defparam \src_data[13]~86 .lut_mask = 16'hFFFE;
defparam \src_data[13]~86 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~87 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_13),
	.datad(out_data_buffer_131),
	.cin(gnd),
	.combout(\src_data[13]~87_combout ),
	.cout());
defparam \src_data[13]~87 .lut_mask = 16'hFFFE;
defparam \src_data[13]~87 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~88 (
	.dataa(\src_data[13]~86_combout ),
	.datab(\src_data[13]~87_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_13),
	.cin(gnd),
	.combout(\src_data[13]~88_combout ),
	.cout());
defparam \src_data[13]~88 .lut_mask = 16'hFFFE;
defparam \src_data[13]~88 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~90 (
	.dataa(src0_valid1),
	.datab(out_valid),
	.datac(out_data_buffer_121),
	.datad(av_readdata_pre_12),
	.cin(gnd),
	.combout(\src_data[12]~90_combout ),
	.cout());
defparam \src_data[12]~90 .lut_mask = 16'hFFFE;
defparam \src_data[12]~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~91 (
	.dataa(read_latency_shift_reg_09),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_121),
	.datad(av_readdata_pre_121),
	.cin(gnd),
	.combout(\src_data[12]~91_combout ),
	.cout());
defparam \src_data[12]~91 .lut_mask = 16'hFFFE;
defparam \src_data[12]~91 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~119 (
	.dataa(out_data_toggle_flopped1),
	.datab(dreg_0),
	.datac(\src_data[12]~91_combout ),
	.datad(out_data_buffer_122),
	.cin(gnd),
	.combout(\src_data[12]~119_combout ),
	.cout());
defparam \src_data[12]~119 .lut_mask = 16'hFFF6;
defparam \src_data[12]~119 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~93 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_111),
	.datad(av_readdata_pre_112),
	.cin(gnd),
	.combout(\src_data[11]~93_combout ),
	.cout());
defparam \src_data[11]~93 .lut_mask = 16'hFFFE;
defparam \src_data[11]~93 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~94 (
	.dataa(\src_data[11]~93_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[11]~94_combout ),
	.cout());
defparam \src_data[11]~94 .lut_mask = 16'hFEFE;
defparam \src_data[11]~94 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~95 (
	.dataa(read_latency_shift_reg_08),
	.datab(read_latency_shift_reg_09),
	.datac(av_readdata_pre_113),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\src_data[11]~95_combout ),
	.cout());
defparam \src_data[11]~95 .lut_mask = 16'hFFFE;
defparam \src_data[11]~95 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~120 (
	.dataa(out_data_toggle_flopped1),
	.datab(dreg_0),
	.datac(\src_data[11]~95_combout ),
	.datad(out_data_buffer_111),
	.cin(gnd),
	.combout(\src_data[11]~120_combout ),
	.cout());
defparam \src_data[11]~120 .lut_mask = 16'hFFF6;
defparam \src_data[11]~120 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~97 (
	.dataa(read_latency_shift_reg_08),
	.datab(read_latency_shift_reg_09),
	.datac(av_readdata_pre_101),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\src_data[10]~97_combout ),
	.cout());
defparam \src_data[10]~97 .lut_mask = 16'hFFFE;
defparam \src_data[10]~97 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~98 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_10),
	.datad(av_readdata_pre_102),
	.cin(gnd),
	.combout(\src_data[10]~98_combout ),
	.cout());
defparam \src_data[10]~98 .lut_mask = 16'hFFFE;
defparam \src_data[10]~98 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~99 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_10),
	.datad(out_data_buffer_101),
	.cin(gnd),
	.combout(\src_data[10]~99_combout ),
	.cout());
defparam \src_data[10]~99 .lut_mask = 16'hFFFE;
defparam \src_data[10]~99 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~100 (
	.dataa(\src_data[10]~98_combout ),
	.datab(\src_data[10]~99_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_10),
	.cin(gnd),
	.combout(\src_data[10]~100_combout ),
	.cout());
defparam \src_data[10]~100 .lut_mask = 16'hFFFE;
defparam \src_data[10]~100 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~102 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_9),
	.datad(av_readdata_pre_91),
	.cin(gnd),
	.combout(\src_data[9]~102_combout ),
	.cout());
defparam \src_data[9]~102 .lut_mask = 16'hFFFE;
defparam \src_data[9]~102 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~103 (
	.dataa(\src_data[9]~102_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_9),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[9]~103_combout ),
	.cout());
defparam \src_data[9]~103 .lut_mask = 16'hFEFE;
defparam \src_data[9]~103 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~104 (
	.dataa(read_latency_shift_reg_06),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_91),
	.datad(readdata_92),
	.cin(gnd),
	.combout(\src_data[9]~104_combout ),
	.cout());
defparam \src_data[9]~104 .lut_mask = 16'hFFFE;
defparam \src_data[9]~104 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~105 (
	.dataa(\src_data[9]~103_combout ),
	.datab(\src_data[9]~104_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_9),
	.cin(gnd),
	.combout(\src_data[9]~105_combout ),
	.cout());
defparam \src_data[9]~105 .lut_mask = 16'hFFFE;
defparam \src_data[9]~105 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~106 (
	.dataa(read_latency_shift_reg_09),
	.datab(out_valid1),
	.datac(out_data_buffer_91),
	.datad(av_readdata_pre_92),
	.cin(gnd),
	.combout(\src_data[9]~106_combout ),
	.cout());
defparam \src_data[9]~106 .lut_mask = 16'hFFFE;
defparam \src_data[9]~106 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~108 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_05),
	.datac(readdata_8),
	.datad(av_readdata_pre_81),
	.cin(gnd),
	.combout(\src_data[8]~108_combout ),
	.cout());
defparam \src_data[8]~108 .lut_mask = 16'hFFFE;
defparam \src_data[8]~108 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~109 (
	.dataa(\src_data[8]~108_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[8]~109_combout ),
	.cout());
defparam \src_data[8]~109 .lut_mask = 16'hFEFE;
defparam \src_data[8]~109 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~110 (
	.dataa(read_latency_shift_reg_06),
	.datab(read_latency_shift_reg_07),
	.datac(readdata_81),
	.datad(readdata_82),
	.cin(gnd),
	.combout(\src_data[8]~110_combout ),
	.cout());
defparam \src_data[8]~110 .lut_mask = 16'hFFFE;
defparam \src_data[8]~110 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~111 (
	.dataa(\src_data[8]~109_combout ),
	.datab(\src_data[8]~110_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_8),
	.cin(gnd),
	.combout(\src_data[8]~111_combout ),
	.cout());
defparam \src_data[8]~111 .lut_mask = 16'hFFFE;
defparam \src_data[8]~111 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~112 (
	.dataa(read_latency_shift_reg_08),
	.datab(read_latency_shift_reg_09),
	.datac(av_readdata_pre_82),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\src_data[8]~112_combout ),
	.cout());
defparam \src_data[8]~112 .lut_mask = 16'hFFFE;
defparam \src_data[8]~112 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~121 (
	.dataa(out_data_toggle_flopped1),
	.datab(dreg_0),
	.datac(\src_data[8]~112_combout ),
	.datad(out_data_buffer_81),
	.cin(gnd),
	.combout(\src_data[8]~121_combout ),
	.cout());
defparam \src_data[8]~121 .lut_mask = 16'hFFF6;
defparam \src_data[8]~121 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_mm_interconnect_0_rsp_mux_001 (
	src1_valid,
	source_addr_1,
	src_payload)/* synthesis synthesis_greybox=1 */;
input 	src1_valid;
input 	source_addr_1;
output 	src_payload;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src_payload~0 (
	.dataa(source_addr_1),
	.datab(src1_valid),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_port_gpio_0 (
	clk,
	W_alu_result_3,
	W_alu_result_2,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	r_sync_rst,
	cp_valid,
	m0_write,
	data,
	d_byteenable_0,
	data1,
	data2,
	data3,
	data4,
	data5,
	data6,
	data7,
	d_byteenable_1,
	data_out_0,
	direction_0,
	data_out_1,
	direction_1,
	data_out_2,
	direction_2,
	data_out_3,
	direction_3,
	data_out_4,
	direction_4,
	data_out_5,
	direction_5,
	data_out_6,
	direction_6,
	data_out_7,
	direction_7,
	data_out_8,
	direction_8,
	data_out_9,
	direction_9,
	data_out_10,
	direction_10,
	data_out_11,
	direction_11,
	data_out_12,
	direction_12,
	data_out_13,
	direction_13,
	data_out_14,
	direction_14,
	data_out_15,
	direction_15,
	data_out_16,
	direction_16,
	data_out_17,
	direction_17,
	data_out_18,
	direction_18,
	data_out_19,
	direction_19,
	data_out_20,
	direction_20,
	data_out_21,
	direction_21,
	data_out_22,
	direction_22,
	data_out_23,
	direction_23,
	data_out_24,
	direction_24,
	data_out_25,
	direction_25,
	data_out_26,
	direction_26,
	data_out_27,
	direction_27,
	data_out_28,
	direction_28,
	data_out_29,
	direction_29,
	data_out_30,
	direction_30,
	data_out_31,
	direction_31,
	d_writedata_10,
	d_byteenable_2,
	d_byteenable_3,
	read_latency_shift_reg,
	d_writedata_8,
	d_writedata_9,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_26,
	readdata_25,
	readdata_24,
	readdata_23,
	readdata_22,
	readdata_21,
	readdata_20,
	readdata_19,
	readdata_18,
	readdata_17,
	readdata_16,
	readdata_15,
	readdata_14,
	readdata_13,
	readdata_12,
	readdata_11,
	readdata_10,
	readdata_9,
	readdata_8,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	port_gpio_0_export_0,
	port_gpio_0_export_1,
	port_gpio_0_export_2,
	port_gpio_0_export_3,
	port_gpio_0_export_4,
	port_gpio_0_export_5,
	port_gpio_0_export_6,
	port_gpio_0_export_7,
	port_gpio_0_export_8,
	port_gpio_0_export_9,
	port_gpio_0_export_10,
	port_gpio_0_export_11,
	port_gpio_0_export_12,
	port_gpio_0_export_13,
	port_gpio_0_export_14,
	port_gpio_0_export_15,
	port_gpio_0_export_16,
	port_gpio_0_export_17,
	port_gpio_0_export_18,
	port_gpio_0_export_19,
	port_gpio_0_export_20,
	port_gpio_0_export_21,
	port_gpio_0_export_22,
	port_gpio_0_export_23,
	port_gpio_0_export_24,
	port_gpio_0_export_25,
	port_gpio_0_export_26,
	port_gpio_0_export_27,
	port_gpio_0_export_28,
	port_gpio_0_export_29,
	port_gpio_0_export_30,
	port_gpio_0_export_31)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	r_sync_rst;
input 	cp_valid;
input 	m0_write;
input 	data;
input 	d_byteenable_0;
input 	data1;
input 	data2;
input 	data3;
input 	data4;
input 	data5;
input 	data6;
input 	data7;
input 	d_byteenable_1;
output 	data_out_0;
output 	direction_0;
output 	data_out_1;
output 	direction_1;
output 	data_out_2;
output 	direction_2;
output 	data_out_3;
output 	direction_3;
output 	data_out_4;
output 	direction_4;
output 	data_out_5;
output 	direction_5;
output 	data_out_6;
output 	direction_6;
output 	data_out_7;
output 	direction_7;
output 	data_out_8;
output 	direction_8;
output 	data_out_9;
output 	direction_9;
output 	data_out_10;
output 	direction_10;
output 	data_out_11;
output 	direction_11;
output 	data_out_12;
output 	direction_12;
output 	data_out_13;
output 	direction_13;
output 	data_out_14;
output 	direction_14;
output 	data_out_15;
output 	direction_15;
output 	data_out_16;
output 	direction_16;
output 	data_out_17;
output 	direction_17;
output 	data_out_18;
output 	direction_18;
output 	data_out_19;
output 	direction_19;
output 	data_out_20;
output 	direction_20;
output 	data_out_21;
output 	direction_21;
output 	data_out_22;
output 	direction_22;
output 	data_out_23;
output 	direction_23;
output 	data_out_24;
output 	direction_24;
output 	data_out_25;
output 	direction_25;
output 	data_out_26;
output 	direction_26;
output 	data_out_27;
output 	direction_27;
output 	data_out_28;
output 	direction_28;
output 	data_out_29;
output 	direction_29;
output 	data_out_30;
output 	direction_30;
output 	data_out_31;
output 	direction_31;
input 	d_writedata_10;
input 	d_byteenable_2;
input 	d_byteenable_3;
input 	read_latency_shift_reg;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_26;
output 	readdata_25;
output 	readdata_24;
output 	readdata_23;
output 	readdata_22;
output 	readdata_21;
output 	readdata_20;
output 	readdata_19;
output 	readdata_18;
output 	readdata_17;
output 	readdata_16;
output 	readdata_15;
output 	readdata_14;
output 	readdata_13;
output 	readdata_12;
output 	readdata_11;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	port_gpio_0_export_0;
input 	port_gpio_0_export_1;
input 	port_gpio_0_export_2;
input 	port_gpio_0_export_3;
input 	port_gpio_0_export_4;
input 	port_gpio_0_export_5;
input 	port_gpio_0_export_6;
input 	port_gpio_0_export_7;
input 	port_gpio_0_export_8;
input 	port_gpio_0_export_9;
input 	port_gpio_0_export_10;
input 	port_gpio_0_export_11;
input 	port_gpio_0_export_12;
input 	port_gpio_0_export_13;
input 	port_gpio_0_export_14;
input 	port_gpio_0_export_15;
input 	port_gpio_0_export_16;
input 	port_gpio_0_export_17;
input 	port_gpio_0_export_18;
input 	port_gpio_0_export_19;
input 	port_gpio_0_export_20;
input 	port_gpio_0_export_21;
input 	port_gpio_0_export_22;
input 	port_gpio_0_export_23;
input 	port_gpio_0_export_24;
input 	port_gpio_0_export_25;
input 	port_gpio_0_export_26;
input 	port_gpio_0_export_27;
input 	port_gpio_0_export_28;
input 	port_gpio_0_export_29;
input 	port_gpio_0_export_30;
input 	port_gpio_0_export_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always2~0_combout ;
wire \data[3]~0_combout ;
wire \data[0]~q ;
wire \always3~0_combout ;
wire \direction~0_combout ;
wire \data[1]~q ;
wire \data[2]~q ;
wire \data[3]~q ;
wire \data[4]~q ;
wire \data[5]~q ;
wire \data[6]~q ;
wire \data[7]~q ;
wire \direction~1_combout ;
wire \data[13]~1_combout ;
wire \data[8]~q ;
wire \direction~2_combout ;
wire \direction~3_combout ;
wire \data[9]~q ;
wire \direction~4_combout ;
wire \data[10]~q ;
wire \direction~5_combout ;
wire \data[11]~q ;
wire \direction~6_combout ;
wire \data[12]~q ;
wire \direction~7_combout ;
wire \data[13]~q ;
wire \direction~8_combout ;
wire \data[14]~q ;
wire \direction~9_combout ;
wire \data[15]~q ;
wire \direction~10_combout ;
wire \data[16]~2_combout ;
wire \data[16]~q ;
wire \direction~11_combout ;
wire \direction~12_combout ;
wire \data[17]~q ;
wire \direction~13_combout ;
wire \data[18]~q ;
wire \direction~14_combout ;
wire \data[19]~q ;
wire \direction~15_combout ;
wire \data[20]~q ;
wire \direction~16_combout ;
wire \data[21]~q ;
wire \direction~17_combout ;
wire \data[22]~q ;
wire \direction~18_combout ;
wire \data[23]~q ;
wire \direction~19_combout ;
wire \data[30]~3_combout ;
wire \data[24]~q ;
wire \direction~20_combout ;
wire \direction~21_combout ;
wire \data[25]~q ;
wire \direction~22_combout ;
wire \data[26]~q ;
wire \direction~23_combout ;
wire \data[27]~q ;
wire \direction~24_combout ;
wire \data[28]~q ;
wire \direction~25_combout ;
wire \data[29]~q ;
wire \direction~26_combout ;
wire \data[30]~q ;
wire \direction~27_combout ;
wire \data[31]~q ;
wire \readdata~0_combout ;
wire \data_in[0]~q ;
wire \readdata~1_combout ;
wire \readdata[10]~2_combout ;
wire \data_in[1]~q ;
wire \readdata~3_combout ;
wire \data_in[2]~q ;
wire \readdata~4_combout ;
wire \data_in[3]~q ;
wire \readdata~5_combout ;
wire \data_in[4]~q ;
wire \readdata~6_combout ;
wire \data_in[5]~q ;
wire \readdata~7_combout ;
wire \data_in[6]~q ;
wire \readdata~8_combout ;
wire \data_in[7]~q ;
wire \readdata~9_combout ;
wire \data_in[26]~q ;
wire \readdata~10_combout ;
wire \data_in[25]~q ;
wire \readdata~11_combout ;
wire \data_in[24]~q ;
wire \readdata~12_combout ;
wire \data_in[23]~q ;
wire \readdata~13_combout ;
wire \data_in[22]~q ;
wire \readdata~14_combout ;
wire \data_in[21]~q ;
wire \readdata~15_combout ;
wire \data_in[20]~q ;
wire \readdata~16_combout ;
wire \data_in[19]~q ;
wire \readdata~17_combout ;
wire \data_in[18]~q ;
wire \readdata~18_combout ;
wire \data_in[17]~q ;
wire \readdata~19_combout ;
wire \data_in[16]~q ;
wire \readdata~20_combout ;
wire \data_in[15]~q ;
wire \readdata~21_combout ;
wire \data_in[14]~q ;
wire \readdata~22_combout ;
wire \data_in[13]~q ;
wire \readdata~23_combout ;
wire \data_in[12]~q ;
wire \readdata~24_combout ;
wire \data_in[11]~q ;
wire \readdata~25_combout ;
wire \data_in[10]~q ;
wire \readdata~26_combout ;
wire \data_in[9]~q ;
wire \readdata~27_combout ;
wire \data_in[8]~q ;
wire \readdata~28_combout ;
wire \data_in[27]~q ;
wire \readdata~29_combout ;
wire \data_in[28]~q ;
wire \readdata~30_combout ;
wire \data_in[29]~q ;
wire \readdata~31_combout ;
wire \data_in[30]~q ;
wire \readdata~32_combout ;
wire \data_in[31]~q ;
wire \readdata~33_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(\data[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \direction[0] (
	.clk(clk),
	.d(data),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~0_combout ),
	.q(direction_0),
	.prn(vcc));
defparam \direction[0] .is_wysiwyg = "true";
defparam \direction[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(\data[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \direction[1] (
	.clk(clk),
	.d(data1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~0_combout ),
	.q(direction_1),
	.prn(vcc));
defparam \direction[1] .is_wysiwyg = "true";
defparam \direction[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(\data[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \direction[2] (
	.clk(clk),
	.d(data2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~0_combout ),
	.q(direction_2),
	.prn(vcc));
defparam \direction[2] .is_wysiwyg = "true";
defparam \direction[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(\data[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \direction[3] (
	.clk(clk),
	.d(data3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~0_combout ),
	.q(direction_3),
	.prn(vcc));
defparam \direction[3] .is_wysiwyg = "true";
defparam \direction[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(\data[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \direction[4] (
	.clk(clk),
	.d(data4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~0_combout ),
	.q(direction_4),
	.prn(vcc));
defparam \direction[4] .is_wysiwyg = "true";
defparam \direction[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(\data[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \direction[5] (
	.clk(clk),
	.d(data5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~0_combout ),
	.q(direction_5),
	.prn(vcc));
defparam \direction[5] .is_wysiwyg = "true";
defparam \direction[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(\data[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \direction[6] (
	.clk(clk),
	.d(data6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~0_combout ),
	.q(direction_6),
	.prn(vcc));
defparam \direction[6] .is_wysiwyg = "true";
defparam \direction[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(\data[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \direction[7] (
	.clk(clk),
	.d(data7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~0_combout ),
	.q(direction_7),
	.prn(vcc));
defparam \direction[7] .is_wysiwyg = "true";
defparam \direction[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(\data[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \direction[8] (
	.clk(clk),
	.d(\direction~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~2_combout ),
	.q(direction_8),
	.prn(vcc));
defparam \direction[8] .is_wysiwyg = "true";
defparam \direction[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(\data[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \direction[9] (
	.clk(clk),
	.d(\direction~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~2_combout ),
	.q(direction_9),
	.prn(vcc));
defparam \direction[9] .is_wysiwyg = "true";
defparam \direction[9] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(\data[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \direction[10] (
	.clk(clk),
	.d(\direction~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~2_combout ),
	.q(direction_10),
	.prn(vcc));
defparam \direction[10] .is_wysiwyg = "true";
defparam \direction[10] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(\data[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \direction[11] (
	.clk(clk),
	.d(\direction~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~2_combout ),
	.q(direction_11),
	.prn(vcc));
defparam \direction[11] .is_wysiwyg = "true";
defparam \direction[11] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk),
	.d(\data[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \direction[12] (
	.clk(clk),
	.d(\direction~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~2_combout ),
	.q(direction_12),
	.prn(vcc));
defparam \direction[12] .is_wysiwyg = "true";
defparam \direction[12] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(\data[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \direction[13] (
	.clk(clk),
	.d(\direction~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~2_combout ),
	.q(direction_13),
	.prn(vcc));
defparam \direction[13] .is_wysiwyg = "true";
defparam \direction[13] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(\data[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \direction[14] (
	.clk(clk),
	.d(\direction~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~2_combout ),
	.q(direction_14),
	.prn(vcc));
defparam \direction[14] .is_wysiwyg = "true";
defparam \direction[14] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(\data[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

dffeas \direction[15] (
	.clk(clk),
	.d(\direction~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~2_combout ),
	.q(direction_15),
	.prn(vcc));
defparam \direction[15] .is_wysiwyg = "true";
defparam \direction[15] .power_up = "low";

dffeas \data_out[16] (
	.clk(clk),
	.d(\data[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_16),
	.prn(vcc));
defparam \data_out[16] .is_wysiwyg = "true";
defparam \data_out[16] .power_up = "low";

dffeas \direction[16] (
	.clk(clk),
	.d(\direction~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~11_combout ),
	.q(direction_16),
	.prn(vcc));
defparam \direction[16] .is_wysiwyg = "true";
defparam \direction[16] .power_up = "low";

dffeas \data_out[17] (
	.clk(clk),
	.d(\data[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_17),
	.prn(vcc));
defparam \data_out[17] .is_wysiwyg = "true";
defparam \data_out[17] .power_up = "low";

dffeas \direction[17] (
	.clk(clk),
	.d(\direction~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~11_combout ),
	.q(direction_17),
	.prn(vcc));
defparam \direction[17] .is_wysiwyg = "true";
defparam \direction[17] .power_up = "low";

dffeas \data_out[18] (
	.clk(clk),
	.d(\data[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_18),
	.prn(vcc));
defparam \data_out[18] .is_wysiwyg = "true";
defparam \data_out[18] .power_up = "low";

dffeas \direction[18] (
	.clk(clk),
	.d(\direction~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~11_combout ),
	.q(direction_18),
	.prn(vcc));
defparam \direction[18] .is_wysiwyg = "true";
defparam \direction[18] .power_up = "low";

dffeas \data_out[19] (
	.clk(clk),
	.d(\data[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_19),
	.prn(vcc));
defparam \data_out[19] .is_wysiwyg = "true";
defparam \data_out[19] .power_up = "low";

dffeas \direction[19] (
	.clk(clk),
	.d(\direction~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~11_combout ),
	.q(direction_19),
	.prn(vcc));
defparam \direction[19] .is_wysiwyg = "true";
defparam \direction[19] .power_up = "low";

dffeas \data_out[20] (
	.clk(clk),
	.d(\data[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_20),
	.prn(vcc));
defparam \data_out[20] .is_wysiwyg = "true";
defparam \data_out[20] .power_up = "low";

dffeas \direction[20] (
	.clk(clk),
	.d(\direction~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~11_combout ),
	.q(direction_20),
	.prn(vcc));
defparam \direction[20] .is_wysiwyg = "true";
defparam \direction[20] .power_up = "low";

dffeas \data_out[21] (
	.clk(clk),
	.d(\data[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_21),
	.prn(vcc));
defparam \data_out[21] .is_wysiwyg = "true";
defparam \data_out[21] .power_up = "low";

dffeas \direction[21] (
	.clk(clk),
	.d(\direction~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~11_combout ),
	.q(direction_21),
	.prn(vcc));
defparam \direction[21] .is_wysiwyg = "true";
defparam \direction[21] .power_up = "low";

dffeas \data_out[22] (
	.clk(clk),
	.d(\data[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_22),
	.prn(vcc));
defparam \data_out[22] .is_wysiwyg = "true";
defparam \data_out[22] .power_up = "low";

dffeas \direction[22] (
	.clk(clk),
	.d(\direction~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~11_combout ),
	.q(direction_22),
	.prn(vcc));
defparam \direction[22] .is_wysiwyg = "true";
defparam \direction[22] .power_up = "low";

dffeas \data_out[23] (
	.clk(clk),
	.d(\data[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_23),
	.prn(vcc));
defparam \data_out[23] .is_wysiwyg = "true";
defparam \data_out[23] .power_up = "low";

dffeas \direction[23] (
	.clk(clk),
	.d(\direction~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~11_combout ),
	.q(direction_23),
	.prn(vcc));
defparam \direction[23] .is_wysiwyg = "true";
defparam \direction[23] .power_up = "low";

dffeas \data_out[24] (
	.clk(clk),
	.d(\data[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_24),
	.prn(vcc));
defparam \data_out[24] .is_wysiwyg = "true";
defparam \data_out[24] .power_up = "low";

dffeas \direction[24] (
	.clk(clk),
	.d(\direction~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~20_combout ),
	.q(direction_24),
	.prn(vcc));
defparam \direction[24] .is_wysiwyg = "true";
defparam \direction[24] .power_up = "low";

dffeas \data_out[25] (
	.clk(clk),
	.d(\data[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_25),
	.prn(vcc));
defparam \data_out[25] .is_wysiwyg = "true";
defparam \data_out[25] .power_up = "low";

dffeas \direction[25] (
	.clk(clk),
	.d(\direction~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~20_combout ),
	.q(direction_25),
	.prn(vcc));
defparam \direction[25] .is_wysiwyg = "true";
defparam \direction[25] .power_up = "low";

dffeas \data_out[26] (
	.clk(clk),
	.d(\data[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_26),
	.prn(vcc));
defparam \data_out[26] .is_wysiwyg = "true";
defparam \data_out[26] .power_up = "low";

dffeas \direction[26] (
	.clk(clk),
	.d(\direction~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~20_combout ),
	.q(direction_26),
	.prn(vcc));
defparam \direction[26] .is_wysiwyg = "true";
defparam \direction[26] .power_up = "low";

dffeas \data_out[27] (
	.clk(clk),
	.d(\data[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_27),
	.prn(vcc));
defparam \data_out[27] .is_wysiwyg = "true";
defparam \data_out[27] .power_up = "low";

dffeas \direction[27] (
	.clk(clk),
	.d(\direction~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~20_combout ),
	.q(direction_27),
	.prn(vcc));
defparam \direction[27] .is_wysiwyg = "true";
defparam \direction[27] .power_up = "low";

dffeas \data_out[28] (
	.clk(clk),
	.d(\data[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_28),
	.prn(vcc));
defparam \data_out[28] .is_wysiwyg = "true";
defparam \data_out[28] .power_up = "low";

dffeas \direction[28] (
	.clk(clk),
	.d(\direction~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~20_combout ),
	.q(direction_28),
	.prn(vcc));
defparam \direction[28] .is_wysiwyg = "true";
defparam \direction[28] .power_up = "low";

dffeas \data_out[29] (
	.clk(clk),
	.d(\data[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_29),
	.prn(vcc));
defparam \data_out[29] .is_wysiwyg = "true";
defparam \data_out[29] .power_up = "low";

dffeas \direction[29] (
	.clk(clk),
	.d(\direction~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~20_combout ),
	.q(direction_29),
	.prn(vcc));
defparam \direction[29] .is_wysiwyg = "true";
defparam \direction[29] .power_up = "low";

dffeas \data_out[30] (
	.clk(clk),
	.d(\data[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_30),
	.prn(vcc));
defparam \data_out[30] .is_wysiwyg = "true";
defparam \data_out[30] .power_up = "low";

dffeas \direction[30] (
	.clk(clk),
	.d(\direction~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~20_combout ),
	.q(direction_30),
	.prn(vcc));
defparam \direction[30] .is_wysiwyg = "true";
defparam \direction[30] .power_up = "low";

dffeas \data_out[31] (
	.clk(clk),
	.d(\data[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_31),
	.prn(vcc));
defparam \data_out[31] .is_wysiwyg = "true";
defparam \data_out[31] .power_up = "low";

dffeas \direction[31] (
	.clk(clk),
	.d(\direction~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\direction~20_combout ),
	.q(direction_31),
	.prn(vcc));
defparam \direction[31] .is_wysiwyg = "true";
defparam \direction[31] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk),
	.d(\readdata~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk),
	.d(\readdata~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk),
	.d(\readdata~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk),
	.d(\readdata~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk),
	.d(\readdata~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk),
	.d(\readdata~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk),
	.d(\readdata~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk),
	.d(\readdata~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk),
	.d(\readdata~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk),
	.d(\readdata~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk),
	.d(\readdata~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk),
	.d(\readdata~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk),
	.d(\readdata~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk),
	.d(\readdata~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk),
	.d(\readdata~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk),
	.d(\readdata~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk),
	.d(\readdata~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk),
	.d(\readdata~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk),
	.d(\readdata~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk),
	.d(\readdata~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk),
	.d(\readdata~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk),
	.d(\readdata~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk),
	.d(\readdata~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk),
	.d(\readdata~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk),
	.d(\readdata~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk),
	.d(\readdata~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk),
	.d(\readdata~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk),
	.d(\readdata~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk),
	.d(\readdata~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk),
	.d(\readdata~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk),
	.d(\readdata~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk),
	.d(\readdata~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[10]~2_combout ),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

cycloneive_lcell_comb \always2~0 (
	.dataa(W_alu_result_3),
	.datab(W_alu_result_2),
	.datac(m0_write),
	.datad(read_latency_shift_reg),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hEFFF;
defparam \always2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data[3]~0 (
	.dataa(\always2~0_combout ),
	.datab(gnd),
	.datac(d_byteenable_0),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data[3]~0_combout ),
	.cout());
defparam \data[3]~0 .lut_mask = 16'hFFF5;
defparam \data[3]~0 .sum_lutc_input = "datac";

dffeas \data[0] (
	.clk(clk),
	.d(data),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[3]~0_combout ),
	.q(\data[0]~q ),
	.prn(vcc));
defparam \data[0] .is_wysiwyg = "true";
defparam \data[0] .power_up = "low";

cycloneive_lcell_comb \always3~0 (
	.dataa(m0_write),
	.datab(W_alu_result_2),
	.datac(read_latency_shift_reg),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\always3~0_combout ),
	.cout());
defparam \always3~0 .lut_mask = 16'hFEFF;
defparam \always3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \direction~0 (
	.dataa(r_sync_rst),
	.datab(d_byteenable_0),
	.datac(\always3~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\direction~0_combout ),
	.cout());
defparam \direction~0 .lut_mask = 16'hFEFE;
defparam \direction~0 .sum_lutc_input = "datac";

dffeas \data[1] (
	.clk(clk),
	.d(data1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[3]~0_combout ),
	.q(\data[1]~q ),
	.prn(vcc));
defparam \data[1] .is_wysiwyg = "true";
defparam \data[1] .power_up = "low";

dffeas \data[2] (
	.clk(clk),
	.d(data2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[3]~0_combout ),
	.q(\data[2]~q ),
	.prn(vcc));
defparam \data[2] .is_wysiwyg = "true";
defparam \data[2] .power_up = "low";

dffeas \data[3] (
	.clk(clk),
	.d(data3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[3]~0_combout ),
	.q(\data[3]~q ),
	.prn(vcc));
defparam \data[3] .is_wysiwyg = "true";
defparam \data[3] .power_up = "low";

dffeas \data[4] (
	.clk(clk),
	.d(data4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[3]~0_combout ),
	.q(\data[4]~q ),
	.prn(vcc));
defparam \data[4] .is_wysiwyg = "true";
defparam \data[4] .power_up = "low";

dffeas \data[5] (
	.clk(clk),
	.d(data5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[3]~0_combout ),
	.q(\data[5]~q ),
	.prn(vcc));
defparam \data[5] .is_wysiwyg = "true";
defparam \data[5] .power_up = "low";

dffeas \data[6] (
	.clk(clk),
	.d(data6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[3]~0_combout ),
	.q(\data[6]~q ),
	.prn(vcc));
defparam \data[6] .is_wysiwyg = "true";
defparam \data[6] .power_up = "low";

dffeas \data[7] (
	.clk(clk),
	.d(data7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[3]~0_combout ),
	.q(\data[7]~q ),
	.prn(vcc));
defparam \data[7] .is_wysiwyg = "true";
defparam \data[7] .power_up = "low";

cycloneive_lcell_comb \direction~1 (
	.dataa(d_writedata_8),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~1_combout ),
	.cout());
defparam \direction~1 .lut_mask = 16'hAAFF;
defparam \direction~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data[13]~1 (
	.dataa(\always2~0_combout ),
	.datab(gnd),
	.datac(d_byteenable_1),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data[13]~1_combout ),
	.cout());
defparam \data[13]~1 .lut_mask = 16'hFFF5;
defparam \data[13]~1 .sum_lutc_input = "datac";

dffeas \data[8] (
	.clk(clk),
	.d(\direction~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[13]~1_combout ),
	.q(\data[8]~q ),
	.prn(vcc));
defparam \data[8] .is_wysiwyg = "true";
defparam \data[8] .power_up = "low";

cycloneive_lcell_comb \direction~2 (
	.dataa(r_sync_rst),
	.datab(d_byteenable_1),
	.datac(\always3~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\direction~2_combout ),
	.cout());
defparam \direction~2 .lut_mask = 16'hFEFE;
defparam \direction~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \direction~3 (
	.dataa(d_writedata_9),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~3_combout ),
	.cout());
defparam \direction~3 .lut_mask = 16'hAAFF;
defparam \direction~3 .sum_lutc_input = "datac";

dffeas \data[9] (
	.clk(clk),
	.d(\direction~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[13]~1_combout ),
	.q(\data[9]~q ),
	.prn(vcc));
defparam \data[9] .is_wysiwyg = "true";
defparam \data[9] .power_up = "low";

cycloneive_lcell_comb \direction~4 (
	.dataa(d_writedata_10),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~4_combout ),
	.cout());
defparam \direction~4 .lut_mask = 16'hAAFF;
defparam \direction~4 .sum_lutc_input = "datac";

dffeas \data[10] (
	.clk(clk),
	.d(\direction~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[13]~1_combout ),
	.q(\data[10]~q ),
	.prn(vcc));
defparam \data[10] .is_wysiwyg = "true";
defparam \data[10] .power_up = "low";

cycloneive_lcell_comb \direction~5 (
	.dataa(d_writedata_11),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~5_combout ),
	.cout());
defparam \direction~5 .lut_mask = 16'hAAFF;
defparam \direction~5 .sum_lutc_input = "datac";

dffeas \data[11] (
	.clk(clk),
	.d(\direction~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[13]~1_combout ),
	.q(\data[11]~q ),
	.prn(vcc));
defparam \data[11] .is_wysiwyg = "true";
defparam \data[11] .power_up = "low";

cycloneive_lcell_comb \direction~6 (
	.dataa(d_writedata_12),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~6_combout ),
	.cout());
defparam \direction~6 .lut_mask = 16'hAAFF;
defparam \direction~6 .sum_lutc_input = "datac";

dffeas \data[12] (
	.clk(clk),
	.d(\direction~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[13]~1_combout ),
	.q(\data[12]~q ),
	.prn(vcc));
defparam \data[12] .is_wysiwyg = "true";
defparam \data[12] .power_up = "low";

cycloneive_lcell_comb \direction~7 (
	.dataa(d_writedata_13),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~7_combout ),
	.cout());
defparam \direction~7 .lut_mask = 16'hAAFF;
defparam \direction~7 .sum_lutc_input = "datac";

dffeas \data[13] (
	.clk(clk),
	.d(\direction~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[13]~1_combout ),
	.q(\data[13]~q ),
	.prn(vcc));
defparam \data[13] .is_wysiwyg = "true";
defparam \data[13] .power_up = "low";

cycloneive_lcell_comb \direction~8 (
	.dataa(d_writedata_14),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~8_combout ),
	.cout());
defparam \direction~8 .lut_mask = 16'hAAFF;
defparam \direction~8 .sum_lutc_input = "datac";

dffeas \data[14] (
	.clk(clk),
	.d(\direction~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[13]~1_combout ),
	.q(\data[14]~q ),
	.prn(vcc));
defparam \data[14] .is_wysiwyg = "true";
defparam \data[14] .power_up = "low";

cycloneive_lcell_comb \direction~9 (
	.dataa(d_writedata_15),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~9_combout ),
	.cout());
defparam \direction~9 .lut_mask = 16'hAAFF;
defparam \direction~9 .sum_lutc_input = "datac";

dffeas \data[15] (
	.clk(clk),
	.d(\direction~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[13]~1_combout ),
	.q(\data[15]~q ),
	.prn(vcc));
defparam \data[15] .is_wysiwyg = "true";
defparam \data[15] .power_up = "low";

cycloneive_lcell_comb \direction~10 (
	.dataa(d_writedata_16),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~10_combout ),
	.cout());
defparam \direction~10 .lut_mask = 16'hAAFF;
defparam \direction~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data[16]~2 (
	.dataa(\always2~0_combout ),
	.datab(gnd),
	.datac(d_byteenable_2),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data[16]~2_combout ),
	.cout());
defparam \data[16]~2 .lut_mask = 16'hFFF5;
defparam \data[16]~2 .sum_lutc_input = "datac";

dffeas \data[16] (
	.clk(clk),
	.d(\direction~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[16]~2_combout ),
	.q(\data[16]~q ),
	.prn(vcc));
defparam \data[16] .is_wysiwyg = "true";
defparam \data[16] .power_up = "low";

cycloneive_lcell_comb \direction~11 (
	.dataa(r_sync_rst),
	.datab(d_byteenable_2),
	.datac(\always3~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\direction~11_combout ),
	.cout());
defparam \direction~11 .lut_mask = 16'hFEFE;
defparam \direction~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \direction~12 (
	.dataa(d_writedata_17),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~12_combout ),
	.cout());
defparam \direction~12 .lut_mask = 16'hAAFF;
defparam \direction~12 .sum_lutc_input = "datac";

dffeas \data[17] (
	.clk(clk),
	.d(\direction~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[16]~2_combout ),
	.q(\data[17]~q ),
	.prn(vcc));
defparam \data[17] .is_wysiwyg = "true";
defparam \data[17] .power_up = "low";

cycloneive_lcell_comb \direction~13 (
	.dataa(d_writedata_18),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~13_combout ),
	.cout());
defparam \direction~13 .lut_mask = 16'hAAFF;
defparam \direction~13 .sum_lutc_input = "datac";

dffeas \data[18] (
	.clk(clk),
	.d(\direction~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[16]~2_combout ),
	.q(\data[18]~q ),
	.prn(vcc));
defparam \data[18] .is_wysiwyg = "true";
defparam \data[18] .power_up = "low";

cycloneive_lcell_comb \direction~14 (
	.dataa(d_writedata_19),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~14_combout ),
	.cout());
defparam \direction~14 .lut_mask = 16'hAAFF;
defparam \direction~14 .sum_lutc_input = "datac";

dffeas \data[19] (
	.clk(clk),
	.d(\direction~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[16]~2_combout ),
	.q(\data[19]~q ),
	.prn(vcc));
defparam \data[19] .is_wysiwyg = "true";
defparam \data[19] .power_up = "low";

cycloneive_lcell_comb \direction~15 (
	.dataa(d_writedata_20),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~15_combout ),
	.cout());
defparam \direction~15 .lut_mask = 16'hAAFF;
defparam \direction~15 .sum_lutc_input = "datac";

dffeas \data[20] (
	.clk(clk),
	.d(\direction~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[16]~2_combout ),
	.q(\data[20]~q ),
	.prn(vcc));
defparam \data[20] .is_wysiwyg = "true";
defparam \data[20] .power_up = "low";

cycloneive_lcell_comb \direction~16 (
	.dataa(d_writedata_21),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~16_combout ),
	.cout());
defparam \direction~16 .lut_mask = 16'hAAFF;
defparam \direction~16 .sum_lutc_input = "datac";

dffeas \data[21] (
	.clk(clk),
	.d(\direction~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[16]~2_combout ),
	.q(\data[21]~q ),
	.prn(vcc));
defparam \data[21] .is_wysiwyg = "true";
defparam \data[21] .power_up = "low";

cycloneive_lcell_comb \direction~17 (
	.dataa(d_writedata_22),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~17_combout ),
	.cout());
defparam \direction~17 .lut_mask = 16'hAAFF;
defparam \direction~17 .sum_lutc_input = "datac";

dffeas \data[22] (
	.clk(clk),
	.d(\direction~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[16]~2_combout ),
	.q(\data[22]~q ),
	.prn(vcc));
defparam \data[22] .is_wysiwyg = "true";
defparam \data[22] .power_up = "low";

cycloneive_lcell_comb \direction~18 (
	.dataa(d_writedata_23),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~18_combout ),
	.cout());
defparam \direction~18 .lut_mask = 16'hAAFF;
defparam \direction~18 .sum_lutc_input = "datac";

dffeas \data[23] (
	.clk(clk),
	.d(\direction~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[16]~2_combout ),
	.q(\data[23]~q ),
	.prn(vcc));
defparam \data[23] .is_wysiwyg = "true";
defparam \data[23] .power_up = "low";

cycloneive_lcell_comb \direction~19 (
	.dataa(d_writedata_24),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~19_combout ),
	.cout());
defparam \direction~19 .lut_mask = 16'hAAFF;
defparam \direction~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data[30]~3 (
	.dataa(\always2~0_combout ),
	.datab(gnd),
	.datac(d_byteenable_3),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data[30]~3_combout ),
	.cout());
defparam \data[30]~3 .lut_mask = 16'hFFF5;
defparam \data[30]~3 .sum_lutc_input = "datac";

dffeas \data[24] (
	.clk(clk),
	.d(\direction~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[30]~3_combout ),
	.q(\data[24]~q ),
	.prn(vcc));
defparam \data[24] .is_wysiwyg = "true";
defparam \data[24] .power_up = "low";

cycloneive_lcell_comb \direction~20 (
	.dataa(r_sync_rst),
	.datab(d_byteenable_3),
	.datac(\always3~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\direction~20_combout ),
	.cout());
defparam \direction~20 .lut_mask = 16'hFEFE;
defparam \direction~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \direction~21 (
	.dataa(d_writedata_25),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~21_combout ),
	.cout());
defparam \direction~21 .lut_mask = 16'hAAFF;
defparam \direction~21 .sum_lutc_input = "datac";

dffeas \data[25] (
	.clk(clk),
	.d(\direction~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[30]~3_combout ),
	.q(\data[25]~q ),
	.prn(vcc));
defparam \data[25] .is_wysiwyg = "true";
defparam \data[25] .power_up = "low";

cycloneive_lcell_comb \direction~22 (
	.dataa(d_writedata_26),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~22_combout ),
	.cout());
defparam \direction~22 .lut_mask = 16'hAAFF;
defparam \direction~22 .sum_lutc_input = "datac";

dffeas \data[26] (
	.clk(clk),
	.d(\direction~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[30]~3_combout ),
	.q(\data[26]~q ),
	.prn(vcc));
defparam \data[26] .is_wysiwyg = "true";
defparam \data[26] .power_up = "low";

cycloneive_lcell_comb \direction~23 (
	.dataa(d_writedata_27),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~23_combout ),
	.cout());
defparam \direction~23 .lut_mask = 16'hAAFF;
defparam \direction~23 .sum_lutc_input = "datac";

dffeas \data[27] (
	.clk(clk),
	.d(\direction~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[30]~3_combout ),
	.q(\data[27]~q ),
	.prn(vcc));
defparam \data[27] .is_wysiwyg = "true";
defparam \data[27] .power_up = "low";

cycloneive_lcell_comb \direction~24 (
	.dataa(d_writedata_28),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~24_combout ),
	.cout());
defparam \direction~24 .lut_mask = 16'hAAFF;
defparam \direction~24 .sum_lutc_input = "datac";

dffeas \data[28] (
	.clk(clk),
	.d(\direction~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[30]~3_combout ),
	.q(\data[28]~q ),
	.prn(vcc));
defparam \data[28] .is_wysiwyg = "true";
defparam \data[28] .power_up = "low";

cycloneive_lcell_comb \direction~25 (
	.dataa(d_writedata_29),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~25_combout ),
	.cout());
defparam \direction~25 .lut_mask = 16'hAAFF;
defparam \direction~25 .sum_lutc_input = "datac";

dffeas \data[29] (
	.clk(clk),
	.d(\direction~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[30]~3_combout ),
	.q(\data[29]~q ),
	.prn(vcc));
defparam \data[29] .is_wysiwyg = "true";
defparam \data[29] .power_up = "low";

cycloneive_lcell_comb \direction~26 (
	.dataa(d_writedata_30),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~26_combout ),
	.cout());
defparam \direction~26 .lut_mask = 16'hAAFF;
defparam \direction~26 .sum_lutc_input = "datac";

dffeas \data[30] (
	.clk(clk),
	.d(\direction~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[30]~3_combout ),
	.q(\data[30]~q ),
	.prn(vcc));
defparam \data[30] .is_wysiwyg = "true";
defparam \data[30] .power_up = "low";

cycloneive_lcell_comb \direction~27 (
	.dataa(d_writedata_31),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\direction~27_combout ),
	.cout());
defparam \direction~27 .lut_mask = 16'hAAFF;
defparam \direction~27 .sum_lutc_input = "datac";

dffeas \data[31] (
	.clk(clk),
	.d(\direction~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[30]~3_combout ),
	.q(\data[31]~q ),
	.prn(vcc));
defparam \data[31] .is_wysiwyg = "true";
defparam \data[31] .power_up = "low";

cycloneive_lcell_comb \readdata~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'h0FFF;
defparam \readdata~0 .sum_lutc_input = "datac";

dffeas \data_in[0] (
	.clk(clk),
	.d(port_gpio_0_export_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[0]~q ),
	.prn(vcc));
defparam \data_in[0] .is_wysiwyg = "true";
defparam \data_in[0] .power_up = "low";

cycloneive_lcell_comb \readdata~1 (
	.dataa(\readdata~0_combout ),
	.datab(direction_0),
	.datac(\data_in[0]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~1_combout ),
	.cout());
defparam \readdata~1 .lut_mask = 16'hFAFC;
defparam \readdata~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[10]~2 (
	.dataa(gnd),
	.datab(cp_valid),
	.datac(read_latency_shift_reg),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata[10]~2_combout ),
	.cout());
defparam \readdata[10]~2 .lut_mask = 16'hFFFC;
defparam \readdata[10]~2 .sum_lutc_input = "datac";

dffeas \data_in[1] (
	.clk(clk),
	.d(port_gpio_0_export_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[1]~q ),
	.prn(vcc));
defparam \data_in[1] .is_wysiwyg = "true";
defparam \data_in[1] .power_up = "low";

cycloneive_lcell_comb \readdata~3 (
	.dataa(\readdata~0_combout ),
	.datab(direction_1),
	.datac(\data_in[1]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hFAFC;
defparam \readdata~3 .sum_lutc_input = "datac";

dffeas \data_in[2] (
	.clk(clk),
	.d(port_gpio_0_export_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[2]~q ),
	.prn(vcc));
defparam \data_in[2] .is_wysiwyg = "true";
defparam \data_in[2] .power_up = "low";

cycloneive_lcell_comb \readdata~4 (
	.dataa(\readdata~0_combout ),
	.datab(direction_2),
	.datac(\data_in[2]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hFAFC;
defparam \readdata~4 .sum_lutc_input = "datac";

dffeas \data_in[3] (
	.clk(clk),
	.d(port_gpio_0_export_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[3]~q ),
	.prn(vcc));
defparam \data_in[3] .is_wysiwyg = "true";
defparam \data_in[3] .power_up = "low";

cycloneive_lcell_comb \readdata~5 (
	.dataa(\readdata~0_combout ),
	.datab(direction_3),
	.datac(\data_in[3]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hFAFC;
defparam \readdata~5 .sum_lutc_input = "datac";

dffeas \data_in[4] (
	.clk(clk),
	.d(port_gpio_0_export_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[4]~q ),
	.prn(vcc));
defparam \data_in[4] .is_wysiwyg = "true";
defparam \data_in[4] .power_up = "low";

cycloneive_lcell_comb \readdata~6 (
	.dataa(\readdata~0_combout ),
	.datab(direction_4),
	.datac(\data_in[4]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hFAFC;
defparam \readdata~6 .sum_lutc_input = "datac";

dffeas \data_in[5] (
	.clk(clk),
	.d(port_gpio_0_export_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[5]~q ),
	.prn(vcc));
defparam \data_in[5] .is_wysiwyg = "true";
defparam \data_in[5] .power_up = "low";

cycloneive_lcell_comb \readdata~7 (
	.dataa(\readdata~0_combout ),
	.datab(direction_5),
	.datac(\data_in[5]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hFAFC;
defparam \readdata~7 .sum_lutc_input = "datac";

dffeas \data_in[6] (
	.clk(clk),
	.d(port_gpio_0_export_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[6]~q ),
	.prn(vcc));
defparam \data_in[6] .is_wysiwyg = "true";
defparam \data_in[6] .power_up = "low";

cycloneive_lcell_comb \readdata~8 (
	.dataa(\readdata~0_combout ),
	.datab(direction_6),
	.datac(\data_in[6]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hFAFC;
defparam \readdata~8 .sum_lutc_input = "datac";

dffeas \data_in[7] (
	.clk(clk),
	.d(port_gpio_0_export_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[7]~q ),
	.prn(vcc));
defparam \data_in[7] .is_wysiwyg = "true";
defparam \data_in[7] .power_up = "low";

cycloneive_lcell_comb \readdata~9 (
	.dataa(\readdata~0_combout ),
	.datab(direction_7),
	.datac(\data_in[7]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~9_combout ),
	.cout());
defparam \readdata~9 .lut_mask = 16'hFAFC;
defparam \readdata~9 .sum_lutc_input = "datac";

dffeas \data_in[26] (
	.clk(clk),
	.d(port_gpio_0_export_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[26]~q ),
	.prn(vcc));
defparam \data_in[26] .is_wysiwyg = "true";
defparam \data_in[26] .power_up = "low";

cycloneive_lcell_comb \readdata~10 (
	.dataa(\readdata~0_combout ),
	.datab(direction_26),
	.datac(\data_in[26]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~10_combout ),
	.cout());
defparam \readdata~10 .lut_mask = 16'hFAFC;
defparam \readdata~10 .sum_lutc_input = "datac";

dffeas \data_in[25] (
	.clk(clk),
	.d(port_gpio_0_export_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[25]~q ),
	.prn(vcc));
defparam \data_in[25] .is_wysiwyg = "true";
defparam \data_in[25] .power_up = "low";

cycloneive_lcell_comb \readdata~11 (
	.dataa(\readdata~0_combout ),
	.datab(direction_25),
	.datac(\data_in[25]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~11_combout ),
	.cout());
defparam \readdata~11 .lut_mask = 16'hFAFC;
defparam \readdata~11 .sum_lutc_input = "datac";

dffeas \data_in[24] (
	.clk(clk),
	.d(port_gpio_0_export_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[24]~q ),
	.prn(vcc));
defparam \data_in[24] .is_wysiwyg = "true";
defparam \data_in[24] .power_up = "low";

cycloneive_lcell_comb \readdata~12 (
	.dataa(\readdata~0_combout ),
	.datab(direction_24),
	.datac(\data_in[24]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~12_combout ),
	.cout());
defparam \readdata~12 .lut_mask = 16'hFAFC;
defparam \readdata~12 .sum_lutc_input = "datac";

dffeas \data_in[23] (
	.clk(clk),
	.d(port_gpio_0_export_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[23]~q ),
	.prn(vcc));
defparam \data_in[23] .is_wysiwyg = "true";
defparam \data_in[23] .power_up = "low";

cycloneive_lcell_comb \readdata~13 (
	.dataa(\readdata~0_combout ),
	.datab(direction_23),
	.datac(\data_in[23]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~13_combout ),
	.cout());
defparam \readdata~13 .lut_mask = 16'hFAFC;
defparam \readdata~13 .sum_lutc_input = "datac";

dffeas \data_in[22] (
	.clk(clk),
	.d(port_gpio_0_export_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[22]~q ),
	.prn(vcc));
defparam \data_in[22] .is_wysiwyg = "true";
defparam \data_in[22] .power_up = "low";

cycloneive_lcell_comb \readdata~14 (
	.dataa(\readdata~0_combout ),
	.datab(direction_22),
	.datac(\data_in[22]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~14_combout ),
	.cout());
defparam \readdata~14 .lut_mask = 16'hFAFC;
defparam \readdata~14 .sum_lutc_input = "datac";

dffeas \data_in[21] (
	.clk(clk),
	.d(port_gpio_0_export_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[21]~q ),
	.prn(vcc));
defparam \data_in[21] .is_wysiwyg = "true";
defparam \data_in[21] .power_up = "low";

cycloneive_lcell_comb \readdata~15 (
	.dataa(\readdata~0_combout ),
	.datab(direction_21),
	.datac(\data_in[21]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~15_combout ),
	.cout());
defparam \readdata~15 .lut_mask = 16'hFAFC;
defparam \readdata~15 .sum_lutc_input = "datac";

dffeas \data_in[20] (
	.clk(clk),
	.d(port_gpio_0_export_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[20]~q ),
	.prn(vcc));
defparam \data_in[20] .is_wysiwyg = "true";
defparam \data_in[20] .power_up = "low";

cycloneive_lcell_comb \readdata~16 (
	.dataa(\readdata~0_combout ),
	.datab(direction_20),
	.datac(\data_in[20]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~16_combout ),
	.cout());
defparam \readdata~16 .lut_mask = 16'hFAFC;
defparam \readdata~16 .sum_lutc_input = "datac";

dffeas \data_in[19] (
	.clk(clk),
	.d(port_gpio_0_export_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[19]~q ),
	.prn(vcc));
defparam \data_in[19] .is_wysiwyg = "true";
defparam \data_in[19] .power_up = "low";

cycloneive_lcell_comb \readdata~17 (
	.dataa(\readdata~0_combout ),
	.datab(direction_19),
	.datac(\data_in[19]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~17_combout ),
	.cout());
defparam \readdata~17 .lut_mask = 16'hFAFC;
defparam \readdata~17 .sum_lutc_input = "datac";

dffeas \data_in[18] (
	.clk(clk),
	.d(port_gpio_0_export_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[18]~q ),
	.prn(vcc));
defparam \data_in[18] .is_wysiwyg = "true";
defparam \data_in[18] .power_up = "low";

cycloneive_lcell_comb \readdata~18 (
	.dataa(\readdata~0_combout ),
	.datab(direction_18),
	.datac(\data_in[18]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~18_combout ),
	.cout());
defparam \readdata~18 .lut_mask = 16'hFAFC;
defparam \readdata~18 .sum_lutc_input = "datac";

dffeas \data_in[17] (
	.clk(clk),
	.d(port_gpio_0_export_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[17]~q ),
	.prn(vcc));
defparam \data_in[17] .is_wysiwyg = "true";
defparam \data_in[17] .power_up = "low";

cycloneive_lcell_comb \readdata~19 (
	.dataa(\readdata~0_combout ),
	.datab(direction_17),
	.datac(\data_in[17]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~19_combout ),
	.cout());
defparam \readdata~19 .lut_mask = 16'hFAFC;
defparam \readdata~19 .sum_lutc_input = "datac";

dffeas \data_in[16] (
	.clk(clk),
	.d(port_gpio_0_export_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[16]~q ),
	.prn(vcc));
defparam \data_in[16] .is_wysiwyg = "true";
defparam \data_in[16] .power_up = "low";

cycloneive_lcell_comb \readdata~20 (
	.dataa(\readdata~0_combout ),
	.datab(direction_16),
	.datac(\data_in[16]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~20_combout ),
	.cout());
defparam \readdata~20 .lut_mask = 16'hFAFC;
defparam \readdata~20 .sum_lutc_input = "datac";

dffeas \data_in[15] (
	.clk(clk),
	.d(port_gpio_0_export_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[15]~q ),
	.prn(vcc));
defparam \data_in[15] .is_wysiwyg = "true";
defparam \data_in[15] .power_up = "low";

cycloneive_lcell_comb \readdata~21 (
	.dataa(\readdata~0_combout ),
	.datab(direction_15),
	.datac(\data_in[15]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~21_combout ),
	.cout());
defparam \readdata~21 .lut_mask = 16'hFAFC;
defparam \readdata~21 .sum_lutc_input = "datac";

dffeas \data_in[14] (
	.clk(clk),
	.d(port_gpio_0_export_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[14]~q ),
	.prn(vcc));
defparam \data_in[14] .is_wysiwyg = "true";
defparam \data_in[14] .power_up = "low";

cycloneive_lcell_comb \readdata~22 (
	.dataa(\readdata~0_combout ),
	.datab(direction_14),
	.datac(\data_in[14]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~22_combout ),
	.cout());
defparam \readdata~22 .lut_mask = 16'hFAFC;
defparam \readdata~22 .sum_lutc_input = "datac";

dffeas \data_in[13] (
	.clk(clk),
	.d(port_gpio_0_export_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[13]~q ),
	.prn(vcc));
defparam \data_in[13] .is_wysiwyg = "true";
defparam \data_in[13] .power_up = "low";

cycloneive_lcell_comb \readdata~23 (
	.dataa(\readdata~0_combout ),
	.datab(direction_13),
	.datac(\data_in[13]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~23_combout ),
	.cout());
defparam \readdata~23 .lut_mask = 16'hFAFC;
defparam \readdata~23 .sum_lutc_input = "datac";

dffeas \data_in[12] (
	.clk(clk),
	.d(port_gpio_0_export_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[12]~q ),
	.prn(vcc));
defparam \data_in[12] .is_wysiwyg = "true";
defparam \data_in[12] .power_up = "low";

cycloneive_lcell_comb \readdata~24 (
	.dataa(\readdata~0_combout ),
	.datab(direction_12),
	.datac(\data_in[12]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~24_combout ),
	.cout());
defparam \readdata~24 .lut_mask = 16'hFAFC;
defparam \readdata~24 .sum_lutc_input = "datac";

dffeas \data_in[11] (
	.clk(clk),
	.d(port_gpio_0_export_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[11]~q ),
	.prn(vcc));
defparam \data_in[11] .is_wysiwyg = "true";
defparam \data_in[11] .power_up = "low";

cycloneive_lcell_comb \readdata~25 (
	.dataa(\readdata~0_combout ),
	.datab(direction_11),
	.datac(\data_in[11]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~25_combout ),
	.cout());
defparam \readdata~25 .lut_mask = 16'hFAFC;
defparam \readdata~25 .sum_lutc_input = "datac";

dffeas \data_in[10] (
	.clk(clk),
	.d(port_gpio_0_export_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[10]~q ),
	.prn(vcc));
defparam \data_in[10] .is_wysiwyg = "true";
defparam \data_in[10] .power_up = "low";

cycloneive_lcell_comb \readdata~26 (
	.dataa(\readdata~0_combout ),
	.datab(direction_10),
	.datac(\data_in[10]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~26_combout ),
	.cout());
defparam \readdata~26 .lut_mask = 16'hFAFC;
defparam \readdata~26 .sum_lutc_input = "datac";

dffeas \data_in[9] (
	.clk(clk),
	.d(port_gpio_0_export_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[9]~q ),
	.prn(vcc));
defparam \data_in[9] .is_wysiwyg = "true";
defparam \data_in[9] .power_up = "low";

cycloneive_lcell_comb \readdata~27 (
	.dataa(\readdata~0_combout ),
	.datab(direction_9),
	.datac(\data_in[9]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~27_combout ),
	.cout());
defparam \readdata~27 .lut_mask = 16'hFAFC;
defparam \readdata~27 .sum_lutc_input = "datac";

dffeas \data_in[8] (
	.clk(clk),
	.d(port_gpio_0_export_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[8]~q ),
	.prn(vcc));
defparam \data_in[8] .is_wysiwyg = "true";
defparam \data_in[8] .power_up = "low";

cycloneive_lcell_comb \readdata~28 (
	.dataa(\readdata~0_combout ),
	.datab(direction_8),
	.datac(\data_in[8]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~28_combout ),
	.cout());
defparam \readdata~28 .lut_mask = 16'hFAFC;
defparam \readdata~28 .sum_lutc_input = "datac";

dffeas \data_in[27] (
	.clk(clk),
	.d(port_gpio_0_export_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[27]~q ),
	.prn(vcc));
defparam \data_in[27] .is_wysiwyg = "true";
defparam \data_in[27] .power_up = "low";

cycloneive_lcell_comb \readdata~29 (
	.dataa(\readdata~0_combout ),
	.datab(direction_27),
	.datac(\data_in[27]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~29_combout ),
	.cout());
defparam \readdata~29 .lut_mask = 16'hFAFC;
defparam \readdata~29 .sum_lutc_input = "datac";

dffeas \data_in[28] (
	.clk(clk),
	.d(port_gpio_0_export_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[28]~q ),
	.prn(vcc));
defparam \data_in[28] .is_wysiwyg = "true";
defparam \data_in[28] .power_up = "low";

cycloneive_lcell_comb \readdata~30 (
	.dataa(\readdata~0_combout ),
	.datab(direction_28),
	.datac(\data_in[28]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~30_combout ),
	.cout());
defparam \readdata~30 .lut_mask = 16'hFAFC;
defparam \readdata~30 .sum_lutc_input = "datac";

dffeas \data_in[29] (
	.clk(clk),
	.d(port_gpio_0_export_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[29]~q ),
	.prn(vcc));
defparam \data_in[29] .is_wysiwyg = "true";
defparam \data_in[29] .power_up = "low";

cycloneive_lcell_comb \readdata~31 (
	.dataa(\readdata~0_combout ),
	.datab(direction_29),
	.datac(\data_in[29]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~31_combout ),
	.cout());
defparam \readdata~31 .lut_mask = 16'hFAFC;
defparam \readdata~31 .sum_lutc_input = "datac";

dffeas \data_in[30] (
	.clk(clk),
	.d(port_gpio_0_export_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[30]~q ),
	.prn(vcc));
defparam \data_in[30] .is_wysiwyg = "true";
defparam \data_in[30] .power_up = "low";

cycloneive_lcell_comb \readdata~32 (
	.dataa(\readdata~0_combout ),
	.datab(direction_30),
	.datac(\data_in[30]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~32_combout ),
	.cout());
defparam \readdata~32 .lut_mask = 16'hFAFC;
defparam \readdata~32 .sum_lutc_input = "datac";

dffeas \data_in[31] (
	.clk(clk),
	.d(port_gpio_0_export_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[31]~q ),
	.prn(vcc));
defparam \data_in[31] .is_wysiwyg = "true";
defparam \data_in[31] .power_up = "low";

cycloneive_lcell_comb \readdata~33 (
	.dataa(\readdata~0_combout ),
	.datab(direction_31),
	.datac(\data_in[31]~q ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~33_combout ),
	.cout());
defparam \readdata~33 .lut_mask = 16'hFAFC;
defparam \readdata~33 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_port_key (
	clk,
	W_alu_result_3,
	W_alu_result_2,
	r_sync_rst,
	cp_valid,
	write,
	readdata_0,
	readdata_1,
	port_key_export_0,
	port_key_export_1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	r_sync_rst;
input 	cp_valid;
input 	write;
output 	readdata_0;
output 	readdata_1;
input 	port_key_export_0;
input 	port_key_export_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_in[0]~0_combout ;
wire \data_in[0]~q ;
wire \readdata~0_combout ;
wire \readdata[0]~1_combout ;
wire \data_in[1]~1_combout ;
wire \data_in[1]~q ;
wire \readdata~2_combout ;


dffeas \readdata[0] (
	.clk(clk),
	.d(\readdata~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

cycloneive_lcell_comb \data_in[0]~0 (
	.dataa(port_key_export_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in[0]~0_combout ),
	.cout());
defparam \data_in[0]~0 .lut_mask = 16'h5555;
defparam \data_in[0]~0 .sum_lutc_input = "datac";

dffeas \data_in[0] (
	.clk(clk),
	.d(\data_in[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[0]~q ),
	.prn(vcc));
defparam \data_in[0] .is_wysiwyg = "true";
defparam \data_in[0] .power_up = "low";

cycloneive_lcell_comb \readdata~0 (
	.dataa(\data_in[0]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hBFFF;
defparam \readdata~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0]~1 (
	.dataa(gnd),
	.datab(cp_valid),
	.datac(write),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata[0]~1_combout ),
	.cout());
defparam \readdata[0]~1 .lut_mask = 16'hFFFC;
defparam \readdata[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in[1]~1 (
	.dataa(port_key_export_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in[1]~1_combout ),
	.cout());
defparam \data_in[1]~1 .lut_mask = 16'h5555;
defparam \data_in[1]~1 .sum_lutc_input = "datac";

dffeas \data_in[1] (
	.clk(clk),
	.d(\data_in[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[1]~q ),
	.prn(vcc));
defparam \data_in[1] .is_wysiwyg = "true";
defparam \data_in[1] .power_up = "low";

cycloneive_lcell_comb \readdata~2 (
	.dataa(\data_in[1]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hBFFF;
defparam \readdata~2 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_port_led (
	clk,
	W_alu_result_3,
	W_alu_result_2,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	r_sync_rst,
	hold_waitrequest,
	d_write,
	write_accepted,
	cp_valid,
	d_writedata_0,
	data,
	d_byteenable_0,
	Equal6,
	read_latency_shift_reg,
	d_writedata_1,
	data1,
	d_writedata_2,
	data2,
	d_writedata_3,
	data3,
	d_writedata_4,
	data4,
	d_writedata_5,
	data5,
	d_writedata_6,
	data6,
	d_writedata_7,
	data7,
	data8,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_3;
input 	W_alu_result_2;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
input 	r_sync_rst;
input 	hold_waitrequest;
input 	d_write;
input 	write_accepted;
input 	cp_valid;
input 	d_writedata_0;
output 	data;
input 	d_byteenable_0;
input 	Equal6;
input 	read_latency_shift_reg;
input 	d_writedata_1;
output 	data1;
input 	d_writedata_2;
output 	data2;
input 	d_writedata_3;
output 	data3;
input 	d_writedata_4;
output 	data4;
input 	d_writedata_5;
output 	data5;
input 	d_writedata_6;
output 	data6;
input 	d_writedata_7;
output 	data7;
output 	data8;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data~1_combout ;
wire \data[6]~2_combout ;
wire \data[0]~q ;
wire \data[1]~q ;
wire \data[2]~q ;
wire \data[3]~q ;
wire \data[4]~q ;
wire \data[5]~q ;
wire \data[6]~q ;
wire \data[7]~q ;
wire \data_in[0]~q ;
wire \readdata~0_combout ;
wire \readdata[0]~1_combout ;
wire \data_in[1]~q ;
wire \readdata~2_combout ;
wire \data_in[2]~q ;
wire \readdata~3_combout ;
wire \data_in[3]~q ;
wire \readdata~4_combout ;
wire \data_in[4]~q ;
wire \readdata~5_combout ;
wire \data_in[5]~q ;
wire \readdata~6_combout ;
wire \data_in[6]~q ;
wire \readdata~7_combout ;
wire \data_in[7]~q ;
wire \readdata~8_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(\data[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(\data[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(\data[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(\data[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(\data[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(\data[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(\data[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(\data[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

cycloneive_lcell_comb \data~0 (
	.dataa(d_writedata_0),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(data),
	.cout());
defparam \data~0 .lut_mask = 16'hAAFF;
defparam \data~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data~3 (
	.dataa(d_writedata_1),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(data1),
	.cout());
defparam \data~3 .lut_mask = 16'hAAFF;
defparam \data~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data~4 (
	.dataa(d_writedata_2),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(data2),
	.cout());
defparam \data~4 .lut_mask = 16'hAAFF;
defparam \data~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data~5 (
	.dataa(d_writedata_3),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(data3),
	.cout());
defparam \data~5 .lut_mask = 16'hAAFF;
defparam \data~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data~6 (
	.dataa(d_writedata_4),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(data4),
	.cout());
defparam \data~6 .lut_mask = 16'hAAFF;
defparam \data~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data~7 (
	.dataa(d_writedata_5),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(data5),
	.cout());
defparam \data~7 .lut_mask = 16'hAAFF;
defparam \data~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data~8 (
	.dataa(d_writedata_6),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(data6),
	.cout());
defparam \data~8 .lut_mask = 16'hAAFF;
defparam \data~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data~9 (
	.dataa(d_writedata_7),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(data7),
	.cout());
defparam \data~9 .lut_mask = 16'hAAFF;
defparam \data~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data~10 (
	.dataa(d_write),
	.datab(d_byteenable_0),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(data8),
	.cout());
defparam \data~10 .lut_mask = 16'hEEFF;
defparam \data~10 .sum_lutc_input = "datac";

dffeas \readdata[0] (
	.clk(clk),
	.d(\readdata~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk),
	.d(\readdata~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk),
	.d(\readdata~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk),
	.d(\readdata~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk),
	.d(\readdata~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk),
	.d(\readdata~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk),
	.d(\readdata~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[0]~1_combout ),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

cycloneive_lcell_comb \data~1 (
	.dataa(write_accepted),
	.datab(hold_waitrequest),
	.datac(d_write),
	.datad(d_byteenable_0),
	.cin(gnd),
	.combout(\data~1_combout ),
	.cout());
defparam \data~1 .lut_mask = 16'hBFFF;
defparam \data~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data[6]~2 (
	.dataa(\data~1_combout ),
	.datab(Equal6),
	.datac(read_latency_shift_reg),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data[6]~2_combout ),
	.cout());
defparam \data[6]~2 .lut_mask = 16'hFFFD;
defparam \data[6]~2 .sum_lutc_input = "datac";

dffeas \data[0] (
	.clk(clk),
	.d(data),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[6]~2_combout ),
	.q(\data[0]~q ),
	.prn(vcc));
defparam \data[0] .is_wysiwyg = "true";
defparam \data[0] .power_up = "low";

dffeas \data[1] (
	.clk(clk),
	.d(data1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[6]~2_combout ),
	.q(\data[1]~q ),
	.prn(vcc));
defparam \data[1] .is_wysiwyg = "true";
defparam \data[1] .power_up = "low";

dffeas \data[2] (
	.clk(clk),
	.d(data2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[6]~2_combout ),
	.q(\data[2]~q ),
	.prn(vcc));
defparam \data[2] .is_wysiwyg = "true";
defparam \data[2] .power_up = "low";

dffeas \data[3] (
	.clk(clk),
	.d(data3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[6]~2_combout ),
	.q(\data[3]~q ),
	.prn(vcc));
defparam \data[3] .is_wysiwyg = "true";
defparam \data[3] .power_up = "low";

dffeas \data[4] (
	.clk(clk),
	.d(data4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[6]~2_combout ),
	.q(\data[4]~q ),
	.prn(vcc));
defparam \data[4] .is_wysiwyg = "true";
defparam \data[4] .power_up = "low";

dffeas \data[5] (
	.clk(clk),
	.d(data5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[6]~2_combout ),
	.q(\data[5]~q ),
	.prn(vcc));
defparam \data[5] .is_wysiwyg = "true";
defparam \data[5] .power_up = "low";

dffeas \data[6] (
	.clk(clk),
	.d(data6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[6]~2_combout ),
	.q(\data[6]~q ),
	.prn(vcc));
defparam \data[6] .is_wysiwyg = "true";
defparam \data[6] .power_up = "low";

dffeas \data[7] (
	.clk(clk),
	.d(data7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data[6]~2_combout ),
	.q(\data[7]~q ),
	.prn(vcc));
defparam \data[7] .is_wysiwyg = "true";
defparam \data[7] .power_up = "low";

dffeas \data_in[0] (
	.clk(clk),
	.d(\data[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[0]~q ),
	.prn(vcc));
defparam \data_in[0] .is_wysiwyg = "true";
defparam \data_in[0] .power_up = "low";

cycloneive_lcell_comb \readdata~0 (
	.dataa(\data_in[0]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hBFFF;
defparam \readdata~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0]~1 (
	.dataa(gnd),
	.datab(cp_valid),
	.datac(read_latency_shift_reg),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata[0]~1_combout ),
	.cout());
defparam \readdata[0]~1 .lut_mask = 16'hFFFC;
defparam \readdata[0]~1 .sum_lutc_input = "datac";

dffeas \data_in[1] (
	.clk(clk),
	.d(\data[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[1]~q ),
	.prn(vcc));
defparam \data_in[1] .is_wysiwyg = "true";
defparam \data_in[1] .power_up = "low";

cycloneive_lcell_comb \readdata~2 (
	.dataa(\data_in[1]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hBFFF;
defparam \readdata~2 .sum_lutc_input = "datac";

dffeas \data_in[2] (
	.clk(clk),
	.d(\data[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[2]~q ),
	.prn(vcc));
defparam \data_in[2] .is_wysiwyg = "true";
defparam \data_in[2] .power_up = "low";

cycloneive_lcell_comb \readdata~3 (
	.dataa(\data_in[2]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hBFFF;
defparam \readdata~3 .sum_lutc_input = "datac";

dffeas \data_in[3] (
	.clk(clk),
	.d(\data[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[3]~q ),
	.prn(vcc));
defparam \data_in[3] .is_wysiwyg = "true";
defparam \data_in[3] .power_up = "low";

cycloneive_lcell_comb \readdata~4 (
	.dataa(\data_in[3]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hBFFF;
defparam \readdata~4 .sum_lutc_input = "datac";

dffeas \data_in[4] (
	.clk(clk),
	.d(\data[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[4]~q ),
	.prn(vcc));
defparam \data_in[4] .is_wysiwyg = "true";
defparam \data_in[4] .power_up = "low";

cycloneive_lcell_comb \readdata~5 (
	.dataa(\data_in[4]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hBFFF;
defparam \readdata~5 .sum_lutc_input = "datac";

dffeas \data_in[5] (
	.clk(clk),
	.d(\data[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[5]~q ),
	.prn(vcc));
defparam \data_in[5] .is_wysiwyg = "true";
defparam \data_in[5] .power_up = "low";

cycloneive_lcell_comb \readdata~6 (
	.dataa(\data_in[5]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hBFFF;
defparam \readdata~6 .sum_lutc_input = "datac";

dffeas \data_in[6] (
	.clk(clk),
	.d(\data[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[6]~q ),
	.prn(vcc));
defparam \data_in[6] .is_wysiwyg = "true";
defparam \data_in[6] .power_up = "low";

cycloneive_lcell_comb \readdata~7 (
	.dataa(\data_in[6]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hBFFF;
defparam \readdata~7 .sum_lutc_input = "datac";

dffeas \data_in[7] (
	.clk(clk),
	.d(\data[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[7]~q ),
	.prn(vcc));
defparam \data_in[7] .is_wysiwyg = "true";
defparam \data_in[7] .power_up = "low";

cycloneive_lcell_comb \readdata~8 (
	.dataa(\data_in[7]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hBFFF;
defparam \readdata~8 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_port_sw (
	clk,
	W_alu_result_3,
	W_alu_result_2,
	r_sync_rst,
	cp_valid,
	write,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	DIP)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	r_sync_rst;
input 	cp_valid;
input 	write;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
input 	[3:0] DIP;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_in[0]~q ;
wire \readdata~0_combout ;
wire \readdata[3]~1_combout ;
wire \data_in[1]~q ;
wire \readdata~2_combout ;
wire \data_in[2]~q ;
wire \readdata~3_combout ;
wire \data_in[3]~q ;
wire \readdata~4_combout ;


dffeas \readdata[0] (
	.clk(clk),
	.d(\readdata~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[3]~1_combout ),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[3]~1_combout ),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk),
	.d(\readdata~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[3]~1_combout ),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk),
	.d(\readdata~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[3]~1_combout ),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \data_in[0] (
	.clk(clk),
	.d(DIP[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[0]~q ),
	.prn(vcc));
defparam \data_in[0] .is_wysiwyg = "true";
defparam \data_in[0] .power_up = "low";

cycloneive_lcell_comb \readdata~0 (
	.dataa(\data_in[0]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hBFFF;
defparam \readdata~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3]~1 (
	.dataa(gnd),
	.datab(cp_valid),
	.datac(write),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata[3]~1_combout ),
	.cout());
defparam \readdata[3]~1 .lut_mask = 16'hFFFC;
defparam \readdata[3]~1 .sum_lutc_input = "datac";

dffeas \data_in[1] (
	.clk(clk),
	.d(DIP[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[1]~q ),
	.prn(vcc));
defparam \data_in[1] .is_wysiwyg = "true";
defparam \data_in[1] .power_up = "low";

cycloneive_lcell_comb \readdata~2 (
	.dataa(\data_in[1]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hBFFF;
defparam \readdata~2 .sum_lutc_input = "datac";

dffeas \data_in[2] (
	.clk(clk),
	.d(DIP[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[2]~q ),
	.prn(vcc));
defparam \data_in[2] .is_wysiwyg = "true";
defparam \data_in[2] .power_up = "low";

cycloneive_lcell_comb \readdata~3 (
	.dataa(\data_in[2]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hBFFF;
defparam \readdata~3 .sum_lutc_input = "datac";

dffeas \data_in[3] (
	.clk(clk),
	.d(DIP[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_in[3]~q ),
	.prn(vcc));
defparam \data_in[3] .is_wysiwyg = "true";
defparam \data_in[3] .power_up = "low";

cycloneive_lcell_comb \readdata~4 (
	.dataa(\data_in[3]~q ),
	.datab(r_sync_rst),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hBFFF;
defparam \readdata~4 .sum_lutc_input = "datac";

endmodule

module niosII_niosII_rs232_0 (
	wire_pll7_clk_0,
	W_alu_result_2,
	readdata_0,
	irq1,
	readdata_1,
	readdata_23,
	readdata_22,
	readdata_21,
	readdata_20,
	readdata_19,
	readdata_18,
	readdata_17,
	readdata_16,
	serial_data_out,
	r_sync_rst,
	d_read,
	read_accepted,
	hold_waitrequest,
	cp_valid,
	data,
	d_byteenable_0,
	Equal9,
	data1,
	data2,
	data3,
	data4,
	data5,
	data6,
	data7,
	Equal12,
	mem_used_1,
	Equal121,
	data_to_uart_0,
	data8,
	read_latency_shift_reg,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	data_to_uart_1,
	readdata_15,
	readdata_9,
	readdata_8,
	data_to_uart_2,
	comb,
	data_to_uart_3,
	data_to_uart_4,
	data_to_uart_5,
	data_to_uart_6,
	data_to_uart_7,
	GND_port,
	rs232_0_RXD)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_2;
output 	readdata_0;
output 	irq1;
output 	readdata_1;
output 	readdata_23;
output 	readdata_22;
output 	readdata_21;
output 	readdata_20;
output 	readdata_19;
output 	readdata_18;
output 	readdata_17;
output 	readdata_16;
output 	serial_data_out;
input 	r_sync_rst;
input 	d_read;
input 	read_accepted;
input 	hold_waitrequest;
input 	cp_valid;
input 	data;
input 	d_byteenable_0;
input 	Equal9;
input 	data1;
input 	data2;
input 	data3;
input 	data4;
input 	data5;
input 	data6;
input 	data7;
input 	Equal12;
input 	mem_used_1;
input 	Equal121;
output 	data_to_uart_0;
input 	data8;
input 	read_latency_shift_reg;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	data_to_uart_1;
output 	readdata_15;
output 	readdata_9;
output 	readdata_8;
output 	data_to_uart_2;
output 	comb;
output 	data_to_uart_3;
output 	data_to_uart_4;
output 	data_to_uart_5;
output 	data_to_uart_6;
output 	data_to_uart_7;
input 	GND_port;
input 	rs232_0_RXD;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write_fifo_write_en~q ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \RS232_Out_Serializer|fifo_write_space[7]~q ;
wire \RS232_Out_Serializer|fifo_write_space[6]~q ;
wire \RS232_Out_Serializer|fifo_write_space[5]~q ;
wire \RS232_Out_Serializer|fifo_write_space[4]~q ;
wire \RS232_Out_Serializer|fifo_write_space[3]~q ;
wire \RS232_Out_Serializer|fifo_write_space[2]~q ;
wire \RS232_Out_Serializer|fifo_write_space[1]~q ;
wire \RS232_Out_Serializer|fifo_write_space[0]~q ;
wire \write_fifo_write_en~0_combout ;
wire \RS232_In_Deserializer|fifo_read_available[7]~q ;
wire \RS232_In_Deserializer|fifo_read_available[6]~q ;
wire \RS232_In_Deserializer|fifo_read_available[5]~q ;
wire \RS232_In_Deserializer|fifo_read_available[4]~q ;
wire \RS232_In_Deserializer|fifo_read_available[3]~q ;
wire \RS232_In_Deserializer|fifo_read_available[2]~q ;
wire \RS232_In_Deserializer|fifo_read_available[1]~q ;
wire \RS232_In_Deserializer|fifo_read_available[0]~q ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \write_fifo_write_en~1_combout ;
wire \write_interrupt_en~0_combout ;
wire \read_interrupt_en~q ;
wire \readdata~0_combout ;
wire \readdata[16]~1_combout ;
wire \read_interrupt~0_combout ;
wire \read_interrupt~q ;
wire \write_interrupt_en~q ;
wire \write_interrupt~0_combout ;
wire \write_interrupt~q ;
wire \irq~0_combout ;
wire \readdata~2_combout ;
wire \readdata~9_combout ;
wire \readdata~10_combout ;
wire \readdata~11_combout ;
wire \readdata~12_combout ;
wire \readdata~13_combout ;
wire \readdata~14_combout ;
wire \readdata~15_combout ;
wire \readdata~16_combout ;
wire \readdata~3_combout ;
wire \readdata~4_combout ;
wire \readdata~5_combout ;
wire \readdata~6_combout ;
wire \readdata~7_combout ;
wire \readdata~8_combout ;
wire \readdata~17_combout ;
wire \readdata~18_combout ;
wire \readdata~19_combout ;


niosII_altera_up_rs232_in_deserializer RS232_In_Deserializer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.W_alu_result_2(W_alu_result_2),
	.q_b_0(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.r_sync_rst(r_sync_rst),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.hold_waitrequest(hold_waitrequest),
	.d_byteenable_0(d_byteenable_0),
	.Equal9(Equal9),
	.mem_used_1(mem_used_1),
	.Equal12(Equal121),
	.fifo_read_available_7(\RS232_In_Deserializer|fifo_read_available[7]~q ),
	.fifo_read_available_6(\RS232_In_Deserializer|fifo_read_available[6]~q ),
	.fifo_read_available_5(\RS232_In_Deserializer|fifo_read_available[5]~q ),
	.fifo_read_available_4(\RS232_In_Deserializer|fifo_read_available[4]~q ),
	.fifo_read_available_3(\RS232_In_Deserializer|fifo_read_available[3]~q ),
	.fifo_read_available_2(\RS232_In_Deserializer|fifo_read_available[2]~q ),
	.fifo_read_available_1(\RS232_In_Deserializer|fifo_read_available[1]~q ),
	.fifo_read_available_0(\RS232_In_Deserializer|fifo_read_available[0]~q ),
	.empty_dff(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.comb(comb),
	.GND_port(GND_port),
	.rs232_0_RXD(rs232_0_RXD));

niosII_altera_up_rs232_out_serializer RS232_Out_Serializer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.write_fifo_write_en(\write_fifo_write_en~q ),
	.fifo_write_space_7(\RS232_Out_Serializer|fifo_write_space[7]~q ),
	.fifo_write_space_6(\RS232_Out_Serializer|fifo_write_space[6]~q ),
	.fifo_write_space_5(\RS232_Out_Serializer|fifo_write_space[5]~q ),
	.fifo_write_space_4(\RS232_Out_Serializer|fifo_write_space[4]~q ),
	.fifo_write_space_3(\RS232_Out_Serializer|fifo_write_space[3]~q ),
	.fifo_write_space_2(\RS232_Out_Serializer|fifo_write_space[2]~q ),
	.fifo_write_space_1(\RS232_Out_Serializer|fifo_write_space[1]~q ),
	.fifo_write_space_0(\RS232_Out_Serializer|fifo_write_space[0]~q ),
	.serial_data_out1(serial_data_out),
	.r_sync_rst(r_sync_rst),
	.data_to_uart_0(data_to_uart_0),
	.data_to_uart_1(data_to_uart_1),
	.data_to_uart_2(data_to_uart_2),
	.data_to_uart_3(data_to_uart_3),
	.data_to_uart_4(data_to_uart_4),
	.data_to_uart_5(data_to_uart_5),
	.data_to_uart_6(data_to_uart_6),
	.data_to_uart_7(data_to_uart_7),
	.GND_port(GND_port));

dffeas write_fifo_write_en(
	.clk(wire_pll7_clk_0),
	.d(\write_fifo_write_en~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\write_fifo_write_en~q ),
	.prn(vcc));
defparam write_fifo_write_en.is_wysiwyg = "true";
defparam write_fifo_write_en.power_up = "low";

cycloneive_lcell_comb \write_fifo_write_en~0 (
	.dataa(cp_valid),
	.datab(data8),
	.datac(read_latency_shift_reg),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\write_fifo_write_en~0_combout ),
	.cout());
defparam \write_fifo_write_en~0 .lut_mask = 16'hFEFF;
defparam \write_fifo_write_en~0 .sum_lutc_input = "datac";

dffeas \readdata[0] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas irq(
	.clk(wire_pll7_clk_0),
	.d(\irq~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(irq1),
	.prn(vcc));
defparam irq.is_wysiwyg = "true";
defparam irq.power_up = "low";

dffeas \readdata[1] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[23] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[22] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[21] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[20] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[19] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[18] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[17] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[16] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \data_to_uart[0] (
	.clk(wire_pll7_clk_0),
	.d(data),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_uart_0),
	.prn(vcc));
defparam \data_to_uart[0] .is_wysiwyg = "true";
defparam \data_to_uart[0] .power_up = "low";

dffeas \readdata[2] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \data_to_uart[1] (
	.clk(wire_pll7_clk_0),
	.d(data1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_uart_1),
	.prn(vcc));
defparam \data_to_uart[1] .is_wysiwyg = "true";
defparam \data_to_uart[1] .power_up = "low";

dffeas \readdata[15] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[9] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[8] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[16]~1_combout ),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \data_to_uart[2] (
	.clk(wire_pll7_clk_0),
	.d(data2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_uart_2),
	.prn(vcc));
defparam \data_to_uart[2] .is_wysiwyg = "true";
defparam \data_to_uart[2] .power_up = "low";

dffeas \data_to_uart[3] (
	.clk(wire_pll7_clk_0),
	.d(data3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_uart_3),
	.prn(vcc));
defparam \data_to_uart[3] .is_wysiwyg = "true";
defparam \data_to_uart[3] .power_up = "low";

dffeas \data_to_uart[4] (
	.clk(wire_pll7_clk_0),
	.d(data4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_uart_4),
	.prn(vcc));
defparam \data_to_uart[4] .is_wysiwyg = "true";
defparam \data_to_uart[4] .power_up = "low";

dffeas \data_to_uart[5] (
	.clk(wire_pll7_clk_0),
	.d(data5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_uart_5),
	.prn(vcc));
defparam \data_to_uart[5] .is_wysiwyg = "true";
defparam \data_to_uart[5] .power_up = "low";

dffeas \data_to_uart[6] (
	.clk(wire_pll7_clk_0),
	.d(data6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_uart_6),
	.prn(vcc));
defparam \data_to_uart[6] .is_wysiwyg = "true";
defparam \data_to_uart[6] .power_up = "low";

dffeas \data_to_uart[7] (
	.clk(wire_pll7_clk_0),
	.d(data7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_to_uart_7),
	.prn(vcc));
defparam \data_to_uart[7] .is_wysiwyg = "true";
defparam \data_to_uart[7] .power_up = "low";

cycloneive_lcell_comb \write_fifo_write_en~1 (
	.dataa(cp_valid),
	.datab(data8),
	.datac(Equal12),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\write_fifo_write_en~1_combout ),
	.cout());
defparam \write_fifo_write_en~1 .lut_mask = 16'hFEFF;
defparam \write_fifo_write_en~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_interrupt_en~0 (
	.dataa(gnd),
	.datab(W_alu_result_2),
	.datac(\write_fifo_write_en~1_combout ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\write_interrupt_en~0_combout ),
	.cout());
defparam \write_interrupt_en~0 .lut_mask = 16'hFFFC;
defparam \write_interrupt_en~0 .sum_lutc_input = "datac";

dffeas read_interrupt_en(
	.clk(wire_pll7_clk_0),
	.d(data),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_interrupt_en~0_combout ),
	.q(\read_interrupt_en~q ),
	.prn(vcc));
defparam read_interrupt_en.is_wysiwyg = "true";
defparam read_interrupt_en.power_up = "low";

cycloneive_lcell_comb \readdata~0 (
	.dataa(\read_interrupt_en~q ),
	.datab(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hAACC;
defparam \readdata~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[16]~1 (
	.dataa(gnd),
	.datab(cp_valid),
	.datac(read_latency_shift_reg),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata[16]~1_combout ),
	.cout());
defparam \readdata[16]~1 .lut_mask = 16'hFFFC;
defparam \readdata[16]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_interrupt~0 (
	.dataa(\read_interrupt_en~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[7]~q ),
	.datac(\RS232_In_Deserializer|fifo_read_available[6]~q ),
	.datad(\RS232_In_Deserializer|fifo_read_available[5]~q ),
	.cin(gnd),
	.combout(\read_interrupt~0_combout ),
	.cout());
defparam \read_interrupt~0 .lut_mask = 16'hFFFE;
defparam \read_interrupt~0 .sum_lutc_input = "datac";

dffeas read_interrupt(
	.clk(wire_pll7_clk_0),
	.d(\read_interrupt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\read_interrupt~q ),
	.prn(vcc));
defparam read_interrupt.is_wysiwyg = "true";
defparam read_interrupt.power_up = "low";

dffeas write_interrupt_en(
	.clk(wire_pll7_clk_0),
	.d(data1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_interrupt_en~0_combout ),
	.q(\write_interrupt_en~q ),
	.prn(vcc));
defparam write_interrupt_en.is_wysiwyg = "true";
defparam write_interrupt_en.power_up = "low";

cycloneive_lcell_comb \write_interrupt~0 (
	.dataa(\write_interrupt_en~q ),
	.datab(\RS232_Out_Serializer|fifo_write_space[7]~q ),
	.datac(\RS232_Out_Serializer|fifo_write_space[6]~q ),
	.datad(\RS232_Out_Serializer|fifo_write_space[5]~q ),
	.cin(gnd),
	.combout(\write_interrupt~0_combout ),
	.cout());
defparam \write_interrupt~0 .lut_mask = 16'hFFFE;
defparam \write_interrupt~0 .sum_lutc_input = "datac";

dffeas write_interrupt(
	.clk(wire_pll7_clk_0),
	.d(\write_interrupt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\write_interrupt~q ),
	.prn(vcc));
defparam write_interrupt.is_wysiwyg = "true";
defparam write_interrupt.power_up = "low";

cycloneive_lcell_comb \irq~0 (
	.dataa(\read_interrupt~q ),
	.datab(\write_interrupt~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\irq~0_combout ),
	.cout());
defparam \irq~0 .lut_mask = 16'hEEEE;
defparam \irq~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~2 (
	.dataa(\write_interrupt_en~q ),
	.datab(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hAACC;
defparam \readdata~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~9 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[7]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[7]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~9_combout ),
	.cout());
defparam \readdata~9 .lut_mask = 16'hAACC;
defparam \readdata~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~10 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[6]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[6]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~10_combout ),
	.cout());
defparam \readdata~10 .lut_mask = 16'hAACC;
defparam \readdata~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~11 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[5]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[5]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~11_combout ),
	.cout());
defparam \readdata~11 .lut_mask = 16'hAACC;
defparam \readdata~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~12 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[4]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[4]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~12_combout ),
	.cout());
defparam \readdata~12 .lut_mask = 16'hAACC;
defparam \readdata~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~13 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[3]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[3]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~13_combout ),
	.cout());
defparam \readdata~13 .lut_mask = 16'hAACC;
defparam \readdata~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~14 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[2]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[2]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~14_combout ),
	.cout());
defparam \readdata~14 .lut_mask = 16'hAACC;
defparam \readdata~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~15 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[1]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[1]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~15_combout ),
	.cout());
defparam \readdata~15 .lut_mask = 16'hAACC;
defparam \readdata~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~16 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[0]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[0]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~16_combout ),
	.cout());
defparam \readdata~16 .lut_mask = 16'hAACC;
defparam \readdata~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~3 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hAFFF;
defparam \readdata~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~4 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hAFFF;
defparam \readdata~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~5 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hAFFF;
defparam \readdata~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~6 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hAFFF;
defparam \readdata~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~7 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hAFFF;
defparam \readdata~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~8 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hAFFF;
defparam \readdata~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~17 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~17_combout ),
	.cout());
defparam \readdata~17 .lut_mask = 16'hAFFF;
defparam \readdata~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~18 (
	.dataa(W_alu_result_2),
	.datab(\write_interrupt~q ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata~18_combout ),
	.cout());
defparam \readdata~18 .lut_mask = 16'hEEFF;
defparam \readdata~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~19 (
	.dataa(W_alu_result_2),
	.datab(\read_interrupt~q ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata~19_combout ),
	.cout());
defparam \readdata~19 .lut_mask = 16'hEEFF;
defparam \readdata~19 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_rs232_in_deserializer (
	wire_pll7_clk_0,
	W_alu_result_2,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	r_sync_rst,
	d_read,
	read_accepted,
	hold_waitrequest,
	d_byteenable_0,
	Equal9,
	mem_used_1,
	Equal12,
	fifo_read_available_7,
	fifo_read_available_6,
	fifo_read_available_5,
	fifo_read_available_4,
	fifo_read_available_3,
	fifo_read_available_2,
	fifo_read_available_1,
	fifo_read_available_0,
	empty_dff,
	comb,
	GND_port,
	rs232_0_RXD)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_2;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	r_sync_rst;
input 	d_read;
input 	read_accepted;
input 	hold_waitrequest;
input 	d_byteenable_0;
input 	Equal9;
input 	mem_used_1;
input 	Equal12;
output 	fifo_read_available_7;
output 	fifo_read_available_6;
output 	fifo_read_available_5;
output 	fifo_read_available_4;
output 	fifo_read_available_3;
output 	fifo_read_available_2;
output 	fifo_read_available_1;
output 	fifo_read_available_0;
output 	empty_dff;
output 	comb;
input 	GND_port;
input 	rs232_0_RXD;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \RS232_In_Counters|baud_clock_falling_edge~q ;
wire \receiving_data~q ;
wire \RS232_In_Counters|all_bits_transmitted~q ;
wire \comb~0_combout ;
wire \data_in_shift_reg[1]~q ;
wire \comb~2_combout ;
wire \comb~3_combout ;
wire \data_in_shift_reg[2]~q ;
wire \data_in_shift_reg[3]~q ;
wire \data_in_shift_reg[4]~q ;
wire \data_in_shift_reg[5]~q ;
wire \data_in_shift_reg[6]~q ;
wire \data_in_shift_reg[7]~q ;
wire \data_in_shift_reg[8]~q ;
wire \data_in_shift_reg~0_combout ;
wire \data_in_shift_reg[6]~1_combout ;
wire \data_in_shift_reg~2_combout ;
wire \data_in_shift_reg~3_combout ;
wire \data_in_shift_reg~4_combout ;
wire \data_in_shift_reg~5_combout ;
wire \data_in_shift_reg~6_combout ;
wire \data_in_shift_reg~7_combout ;
wire \data_in_shift_reg[9]~q ;
wire \data_in_shift_reg~8_combout ;
wire \data_in_shift_reg~9_combout ;
wire \receiving_data~0_combout ;
wire \fifo_read_available~0_combout ;
wire \fifo_read_available~1_combout ;
wire \fifo_read_available~2_combout ;
wire \fifo_read_available~3_combout ;
wire \fifo_read_available~4_combout ;
wire \fifo_read_available~5_combout ;
wire \fifo_read_available~6_combout ;
wire \fifo_read_available~7_combout ;


niosII_altera_up_sync_fifo RS232_In_FIFO(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.full_dff(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.counter_reg_bit_6(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.counter_reg_bit_5(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.all_bits_transmitted(\RS232_In_Counters|all_bits_transmitted~q ),
	.comb(\comb~0_combout ),
	.data_in_shift_reg_1(\data_in_shift_reg[1]~q ),
	.comb1(\comb~3_combout ),
	.data_in_shift_reg_2(\data_in_shift_reg[2]~q ),
	.data_in_shift_reg_3(\data_in_shift_reg[3]~q ),
	.data_in_shift_reg_4(\data_in_shift_reg[4]~q ),
	.data_in_shift_reg_5(\data_in_shift_reg[5]~q ),
	.data_in_shift_reg_6(\data_in_shift_reg[6]~q ),
	.data_in_shift_reg_7(\data_in_shift_reg[7]~q ),
	.data_in_shift_reg_8(\data_in_shift_reg[8]~q ),
	.GND_port(GND_port));

niosII_altera_up_rs232_counters RS232_In_Counters(
	.clk(wire_pll7_clk_0),
	.baud_clock_falling_edge1(\RS232_In_Counters|baud_clock_falling_edge~q ),
	.receiving_data(\receiving_data~q ),
	.r_sync_rst(r_sync_rst),
	.all_bits_transmitted1(\RS232_In_Counters|all_bits_transmitted~q ));

dffeas receiving_data(
	.clk(wire_pll7_clk_0),
	.d(\receiving_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\receiving_data~q ),
	.prn(vcc));
defparam receiving_data.is_wysiwyg = "true";
defparam receiving_data.power_up = "low";

cycloneive_lcell_comb \comb~0 (
	.dataa(\RS232_In_Counters|all_bits_transmitted~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hAAFF;
defparam \comb~0 .sum_lutc_input = "datac";

dffeas \data_in_shift_reg[1] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[6]~1_combout ),
	.q(\data_in_shift_reg[1]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[1] .is_wysiwyg = "true";
defparam \data_in_shift_reg[1] .power_up = "low";

cycloneive_lcell_comb \comb~2 (
	.dataa(empty_dff),
	.datab(comb),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\comb~2_combout ),
	.cout());
defparam \comb~2 .lut_mask = 16'hEEFF;
defparam \comb~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~3 (
	.dataa(Equal9),
	.datab(Equal12),
	.datac(\comb~2_combout ),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\comb~3_combout ),
	.cout());
defparam \comb~3 .lut_mask = 16'hFEFF;
defparam \comb~3 .sum_lutc_input = "datac";

dffeas \data_in_shift_reg[2] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[6]~1_combout ),
	.q(\data_in_shift_reg[2]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[2] .is_wysiwyg = "true";
defparam \data_in_shift_reg[2] .power_up = "low";

dffeas \data_in_shift_reg[3] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[6]~1_combout ),
	.q(\data_in_shift_reg[3]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[3] .is_wysiwyg = "true";
defparam \data_in_shift_reg[3] .power_up = "low";

dffeas \data_in_shift_reg[4] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[6]~1_combout ),
	.q(\data_in_shift_reg[4]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[4] .is_wysiwyg = "true";
defparam \data_in_shift_reg[4] .power_up = "low";

dffeas \data_in_shift_reg[5] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[6]~1_combout ),
	.q(\data_in_shift_reg[5]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[5] .is_wysiwyg = "true";
defparam \data_in_shift_reg[5] .power_up = "low";

dffeas \data_in_shift_reg[6] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[6]~1_combout ),
	.q(\data_in_shift_reg[6]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[6] .is_wysiwyg = "true";
defparam \data_in_shift_reg[6] .power_up = "low";

dffeas \data_in_shift_reg[7] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[6]~1_combout ),
	.q(\data_in_shift_reg[7]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[7] .is_wysiwyg = "true";
defparam \data_in_shift_reg[7] .power_up = "low";

dffeas \data_in_shift_reg[8] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[6]~1_combout ),
	.q(\data_in_shift_reg[8]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[8] .is_wysiwyg = "true";
defparam \data_in_shift_reg[8] .power_up = "low";

cycloneive_lcell_comb \data_in_shift_reg~0 (
	.dataa(\data_in_shift_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~0_combout ),
	.cout());
defparam \data_in_shift_reg~0 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg[6]~1 (
	.dataa(r_sync_rst),
	.datab(\RS232_In_Counters|baud_clock_falling_edge~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_shift_reg[6]~1_combout ),
	.cout());
defparam \data_in_shift_reg[6]~1 .lut_mask = 16'hEEEE;
defparam \data_in_shift_reg[6]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~2 (
	.dataa(\data_in_shift_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~2_combout ),
	.cout());
defparam \data_in_shift_reg~2 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~3 (
	.dataa(\data_in_shift_reg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~3_combout ),
	.cout());
defparam \data_in_shift_reg~3 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~4 (
	.dataa(\data_in_shift_reg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~4_combout ),
	.cout());
defparam \data_in_shift_reg~4 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~5 (
	.dataa(\data_in_shift_reg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~5_combout ),
	.cout());
defparam \data_in_shift_reg~5 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~6 (
	.dataa(\data_in_shift_reg[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~6_combout ),
	.cout());
defparam \data_in_shift_reg~6 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~7 (
	.dataa(\data_in_shift_reg[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~7_combout ),
	.cout());
defparam \data_in_shift_reg~7 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~7 .sum_lutc_input = "datac";

dffeas \data_in_shift_reg[9] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[6]~1_combout ),
	.q(\data_in_shift_reg[9]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[9] .is_wysiwyg = "true";
defparam \data_in_shift_reg[9] .power_up = "low";

cycloneive_lcell_comb \data_in_shift_reg~8 (
	.dataa(\data_in_shift_reg[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~8_combout ),
	.cout());
defparam \data_in_shift_reg~8 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~9 (
	.dataa(rs232_0_RXD),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~9_combout ),
	.cout());
defparam \data_in_shift_reg~9 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \receiving_data~0 (
	.dataa(\receiving_data~q ),
	.datab(gnd),
	.datac(rs232_0_RXD),
	.datad(\RS232_In_Counters|all_bits_transmitted~q ),
	.cin(gnd),
	.combout(\receiving_data~0_combout ),
	.cout());
defparam \receiving_data~0 .lut_mask = 16'hAFFF;
defparam \receiving_data~0 .sum_lutc_input = "datac";

dffeas \fifo_read_available[7] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_7),
	.prn(vcc));
defparam \fifo_read_available[7] .is_wysiwyg = "true";
defparam \fifo_read_available[7] .power_up = "low";

dffeas \fifo_read_available[6] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_6),
	.prn(vcc));
defparam \fifo_read_available[6] .is_wysiwyg = "true";
defparam \fifo_read_available[6] .power_up = "low";

dffeas \fifo_read_available[5] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_5),
	.prn(vcc));
defparam \fifo_read_available[5] .is_wysiwyg = "true";
defparam \fifo_read_available[5] .power_up = "low";

dffeas \fifo_read_available[4] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_4),
	.prn(vcc));
defparam \fifo_read_available[4] .is_wysiwyg = "true";
defparam \fifo_read_available[4] .power_up = "low";

dffeas \fifo_read_available[3] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_3),
	.prn(vcc));
defparam \fifo_read_available[3] .is_wysiwyg = "true";
defparam \fifo_read_available[3] .power_up = "low";

dffeas \fifo_read_available[2] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_2),
	.prn(vcc));
defparam \fifo_read_available[2] .is_wysiwyg = "true";
defparam \fifo_read_available[2] .power_up = "low";

dffeas \fifo_read_available[1] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_1),
	.prn(vcc));
defparam \fifo_read_available[1] .is_wysiwyg = "true";
defparam \fifo_read_available[1] .power_up = "low";

dffeas \fifo_read_available[0] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_0),
	.prn(vcc));
defparam \fifo_read_available[0] .is_wysiwyg = "true";
defparam \fifo_read_available[0] .power_up = "low";

cycloneive_lcell_comb \comb~1 (
	.dataa(hold_waitrequest),
	.datab(d_read),
	.datac(d_byteenable_0),
	.datad(read_accepted),
	.cin(gnd),
	.combout(comb),
	.cout());
defparam \comb~1 .lut_mask = 16'hFEFF;
defparam \comb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~0 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~0_combout ),
	.cout());
defparam \fifo_read_available~0 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~1 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~1_combout ),
	.cout());
defparam \fifo_read_available~1 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~2 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~2_combout ),
	.cout());
defparam \fifo_read_available~2 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~3 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~3_combout ),
	.cout());
defparam \fifo_read_available~3 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~4 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~4_combout ),
	.cout());
defparam \fifo_read_available~4 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~5 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~5_combout ),
	.cout());
defparam \fifo_read_available~5 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~6 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~6_combout ),
	.cout());
defparam \fifo_read_available~6 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~7 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~7_combout ),
	.cout());
defparam \fifo_read_available~7 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~7 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_rs232_counters (
	clk,
	baud_clock_falling_edge1,
	receiving_data,
	r_sync_rst,
	all_bits_transmitted1)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	baud_clock_falling_edge1;
input 	receiving_data;
input 	r_sync_rst;
output 	all_bits_transmitted1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \baud_counter[0]~10_combout ;
wire \baud_counter[5]~22 ;
wire \baud_counter[6]~23_combout ;
wire \baud_counter[6]~q ;
wire \Equal0~0_combout ;
wire \baud_counter[6]~24 ;
wire \baud_counter[7]~25_combout ;
wire \baud_counter[7]~q ;
wire \baud_counter[7]~26 ;
wire \baud_counter[8]~27_combout ;
wire \baud_counter[8]~q ;
wire \baud_counter[8]~28 ;
wire \baud_counter[9]~29_combout ;
wire \baud_counter[9]~q ;
wire \Equal0~1_combout ;
wire \baud_counter[8]~14_combout ;
wire \baud_counter[0]~q ;
wire \baud_counter[0]~11 ;
wire \baud_counter[1]~12_combout ;
wire \baud_counter[1]~q ;
wire \baud_counter[1]~13 ;
wire \baud_counter[2]~15_combout ;
wire \baud_counter[2]~q ;
wire \baud_counter[2]~16 ;
wire \baud_counter[3]~17_combout ;
wire \baud_counter[3]~q ;
wire \baud_counter[3]~18 ;
wire \baud_counter[4]~19_combout ;
wire \baud_counter[4]~q ;
wire \baud_counter[4]~20 ;
wire \baud_counter[5]~21_combout ;
wire \baud_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \Equal1~2_combout ;
wire \bit_counter[2]~0_combout ;
wire \bit_counter[0]~2_combout ;
wire \bit_counter[0]~q ;
wire \bit_counter[1]~3_combout ;
wire \bit_counter[1]~q ;
wire \Add1~0_combout ;
wire \bit_counter[2]~1_combout ;
wire \bit_counter[2]~q ;
wire \Add1~1_combout ;
wire \bit_counter[3]~4_combout ;
wire \bit_counter[3]~q ;
wire \Equal2~0_combout ;
wire \all_bits_transmitted~0_combout ;


dffeas baud_clock_falling_edge(
	.clk(clk),
	.d(\Equal1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(baud_clock_falling_edge1),
	.prn(vcc));
defparam baud_clock_falling_edge.is_wysiwyg = "true";
defparam baud_clock_falling_edge.power_up = "low";

dffeas all_bits_transmitted(
	.clk(clk),
	.d(\all_bits_transmitted~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(all_bits_transmitted1),
	.prn(vcc));
defparam all_bits_transmitted.is_wysiwyg = "true";
defparam all_bits_transmitted.power_up = "low";

cycloneive_lcell_comb \baud_counter[0]~10 (
	.dataa(\baud_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\baud_counter[0]~10_combout ),
	.cout(\baud_counter[0]~11 ));
defparam \baud_counter[0]~10 .lut_mask = 16'h55AA;
defparam \baud_counter[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[5]~21 (
	.dataa(\baud_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[4]~20 ),
	.combout(\baud_counter[5]~21_combout ),
	.cout(\baud_counter[5]~22 ));
defparam \baud_counter[5]~21 .lut_mask = 16'h5A5F;
defparam \baud_counter[5]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \baud_counter[6]~23 (
	.dataa(\baud_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[5]~22 ),
	.combout(\baud_counter[6]~23_combout ),
	.cout(\baud_counter[6]~24 ));
defparam \baud_counter[6]~23 .lut_mask = 16'h5AAF;
defparam \baud_counter[6]~23 .sum_lutc_input = "cin";

dffeas \baud_counter[6] (
	.clk(clk),
	.d(\baud_counter[6]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[6]~q ),
	.prn(vcc));
defparam \baud_counter[6] .is_wysiwyg = "true";
defparam \baud_counter[6] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\baud_counter[1]~q ),
	.datab(\baud_counter[4]~q ),
	.datac(\baud_counter[2]~q ),
	.datad(\baud_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[7]~25 (
	.dataa(\baud_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[6]~24 ),
	.combout(\baud_counter[7]~25_combout ),
	.cout(\baud_counter[7]~26 ));
defparam \baud_counter[7]~25 .lut_mask = 16'h5A5F;
defparam \baud_counter[7]~25 .sum_lutc_input = "cin";

dffeas \baud_counter[7] (
	.clk(clk),
	.d(\baud_counter[7]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[7]~q ),
	.prn(vcc));
defparam \baud_counter[7] .is_wysiwyg = "true";
defparam \baud_counter[7] .power_up = "low";

cycloneive_lcell_comb \baud_counter[8]~27 (
	.dataa(\baud_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[7]~26 ),
	.combout(\baud_counter[8]~27_combout ),
	.cout(\baud_counter[8]~28 ));
defparam \baud_counter[8]~27 .lut_mask = 16'h5AAF;
defparam \baud_counter[8]~27 .sum_lutc_input = "cin";

dffeas \baud_counter[8] (
	.clk(clk),
	.d(\baud_counter[8]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[8]~q ),
	.prn(vcc));
defparam \baud_counter[8] .is_wysiwyg = "true";
defparam \baud_counter[8] .power_up = "low";

cycloneive_lcell_comb \baud_counter[9]~29 (
	.dataa(\baud_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\baud_counter[8]~28 ),
	.combout(\baud_counter[9]~29_combout ),
	.cout());
defparam \baud_counter[9]~29 .lut_mask = 16'h5A5A;
defparam \baud_counter[9]~29 .sum_lutc_input = "cin";

dffeas \baud_counter[9] (
	.clk(clk),
	.d(\baud_counter[9]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[9]~q ),
	.prn(vcc));
defparam \baud_counter[9] .is_wysiwyg = "true";
defparam \baud_counter[9] .power_up = "low";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\Equal0~0_combout ),
	.datab(\baud_counter[7]~q ),
	.datac(\Equal1~0_combout ),
	.datad(\baud_counter[9]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[8]~14 (
	.dataa(\Equal0~1_combout ),
	.datab(receiving_data),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\baud_counter[8]~14_combout ),
	.cout());
defparam \baud_counter[8]~14 .lut_mask = 16'hFF77;
defparam \baud_counter[8]~14 .sum_lutc_input = "datac";

dffeas \baud_counter[0] (
	.clk(clk),
	.d(\baud_counter[0]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[0]~q ),
	.prn(vcc));
defparam \baud_counter[0] .is_wysiwyg = "true";
defparam \baud_counter[0] .power_up = "low";

cycloneive_lcell_comb \baud_counter[1]~12 (
	.dataa(\baud_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[0]~11 ),
	.combout(\baud_counter[1]~12_combout ),
	.cout(\baud_counter[1]~13 ));
defparam \baud_counter[1]~12 .lut_mask = 16'h5A5F;
defparam \baud_counter[1]~12 .sum_lutc_input = "cin";

dffeas \baud_counter[1] (
	.clk(clk),
	.d(\baud_counter[1]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[1]~q ),
	.prn(vcc));
defparam \baud_counter[1] .is_wysiwyg = "true";
defparam \baud_counter[1] .power_up = "low";

cycloneive_lcell_comb \baud_counter[2]~15 (
	.dataa(\baud_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[1]~13 ),
	.combout(\baud_counter[2]~15_combout ),
	.cout(\baud_counter[2]~16 ));
defparam \baud_counter[2]~15 .lut_mask = 16'h5AAF;
defparam \baud_counter[2]~15 .sum_lutc_input = "cin";

dffeas \baud_counter[2] (
	.clk(clk),
	.d(\baud_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[2]~q ),
	.prn(vcc));
defparam \baud_counter[2] .is_wysiwyg = "true";
defparam \baud_counter[2] .power_up = "low";

cycloneive_lcell_comb \baud_counter[3]~17 (
	.dataa(\baud_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[2]~16 ),
	.combout(\baud_counter[3]~17_combout ),
	.cout(\baud_counter[3]~18 ));
defparam \baud_counter[3]~17 .lut_mask = 16'h5A5F;
defparam \baud_counter[3]~17 .sum_lutc_input = "cin";

dffeas \baud_counter[3] (
	.clk(clk),
	.d(\baud_counter[3]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[3]~q ),
	.prn(vcc));
defparam \baud_counter[3] .is_wysiwyg = "true";
defparam \baud_counter[3] .power_up = "low";

cycloneive_lcell_comb \baud_counter[4]~19 (
	.dataa(\baud_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[3]~18 ),
	.combout(\baud_counter[4]~19_combout ),
	.cout(\baud_counter[4]~20 ));
defparam \baud_counter[4]~19 .lut_mask = 16'h5AAF;
defparam \baud_counter[4]~19 .sum_lutc_input = "cin";

dffeas \baud_counter[4] (
	.clk(clk),
	.d(\baud_counter[4]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[4]~q ),
	.prn(vcc));
defparam \baud_counter[4] .is_wysiwyg = "true";
defparam \baud_counter[4] .power_up = "low";

dffeas \baud_counter[5] (
	.clk(clk),
	.d(\baud_counter[5]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[8]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[5]~q ),
	.prn(vcc));
defparam \baud_counter[5] .is_wysiwyg = "true";
defparam \baud_counter[5] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\baud_counter[5]~q ),
	.datab(\baud_counter[8]~q ),
	.datac(\baud_counter[0]~q ),
	.datad(\baud_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(\baud_counter[1]~q ),
	.datab(\baud_counter[4]~q ),
	.datac(\baud_counter[2]~q ),
	.datad(\baud_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hEFFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(\Equal1~0_combout ),
	.datab(\baud_counter[7]~q ),
	.datac(\Equal1~1_combout ),
	.datad(\baud_counter[9]~q ),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'hFEFF;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[2]~0 (
	.dataa(\Equal2~0_combout ),
	.datab(receiving_data),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\bit_counter[2]~0_combout ),
	.cout());
defparam \bit_counter[2]~0 .lut_mask = 16'hEEFF;
defparam \bit_counter[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[0]~2 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[0]~q ),
	.datac(\Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\bit_counter[0]~2_combout ),
	.cout());
defparam \bit_counter[0]~2 .lut_mask = 16'hBEBE;
defparam \bit_counter[0]~2 .sum_lutc_input = "datac";

dffeas \bit_counter[0] (
	.clk(clk),
	.d(\bit_counter[0]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[0]~q ),
	.prn(vcc));
defparam \bit_counter[0] .is_wysiwyg = "true";
defparam \bit_counter[0] .power_up = "low";

cycloneive_lcell_comb \bit_counter[1]~3 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[1]~q ),
	.datac(\Equal0~1_combout ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\bit_counter[1]~3_combout ),
	.cout());
defparam \bit_counter[1]~3 .lut_mask = 16'hEBBE;
defparam \bit_counter[1]~3 .sum_lutc_input = "datac";

dffeas \bit_counter[1] (
	.clk(clk),
	.d(\bit_counter[1]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[1]~q ),
	.prn(vcc));
defparam \bit_counter[1] .is_wysiwyg = "true";
defparam \bit_counter[1] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(\bit_counter[2]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'hC33C;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[2]~1 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[2]~q ),
	.datac(\Add1~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\bit_counter[2]~1_combout ),
	.cout());
defparam \bit_counter[2]~1 .lut_mask = 16'hFAFC;
defparam \bit_counter[2]~1 .sum_lutc_input = "datac";

dffeas \bit_counter[2] (
	.clk(clk),
	.d(\bit_counter[2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[2]~q ),
	.prn(vcc));
defparam \bit_counter[2] .is_wysiwyg = "true";
defparam \bit_counter[2] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(\bit_counter[3]~q ),
	.datab(\bit_counter[2]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[3]~4 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[3]~q ),
	.datac(\Add1~1_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\bit_counter[3]~4_combout ),
	.cout());
defparam \bit_counter[3]~4 .lut_mask = 16'hFAFC;
defparam \bit_counter[3]~4 .sum_lutc_input = "datac";

dffeas \bit_counter[3] (
	.clk(clk),
	.d(\bit_counter[3]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[3]~q ),
	.prn(vcc));
defparam \bit_counter[3] .is_wysiwyg = "true";
defparam \bit_counter[3] .power_up = "low";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(\bit_counter[2]~q ),
	.datab(\bit_counter[0]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hEFFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \all_bits_transmitted~0 (
	.dataa(r_sync_rst),
	.datab(\Equal2~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\all_bits_transmitted~0_combout ),
	.cout());
defparam \all_bits_transmitted~0 .lut_mask = 16'h7777;
defparam \all_bits_transmitted~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_sync_fifo (
	wire_pll7_clk_0,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	full_dff,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	empty_dff,
	all_bits_transmitted,
	comb,
	data_in_shift_reg_1,
	comb1,
	data_in_shift_reg_2,
	data_in_shift_reg_3,
	data_in_shift_reg_4,
	data_in_shift_reg_5,
	data_in_shift_reg_6,
	data_in_shift_reg_7,
	data_in_shift_reg_8,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	full_dff;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
output 	empty_dff;
input 	all_bits_transmitted;
input 	comb;
input 	data_in_shift_reg_1;
input 	comb1;
input 	data_in_shift_reg_2;
input 	data_in_shift_reg_3;
input 	data_in_shift_reg_4;
input 	data_in_shift_reg_5;
input 	data_in_shift_reg_6;
input 	data_in_shift_reg_7;
input 	data_in_shift_reg_8;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_3 Sync_FIFO(
	.clock(wire_pll7_clk_0),
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.full_dff(full_dff),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.all_bits_transmitted(all_bits_transmitted),
	.wrreq(comb),
	.data({data_in_shift_reg_8,data_in_shift_reg_7,data_in_shift_reg_6,data_in_shift_reg_5,data_in_shift_reg_4,data_in_shift_reg_3,data_in_shift_reg_2,data_in_shift_reg_1}),
	.comb(comb1),
	.GND_port(GND_port));

endmodule

module niosII_scfifo_3 (
	clock,
	q,
	full_dff,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	empty_dff,
	all_bits_transmitted,
	wrreq,
	data,
	comb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
output 	full_dff;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
output 	empty_dff;
input 	all_bits_transmitted;
input 	wrreq;
input 	[7:0] data;
input 	comb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_a341 auto_generated(
	.clock(clock),
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.full_dff(full_dff),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.all_bits_transmitted(all_bits_transmitted),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.comb(comb),
	.GND_port(GND_port));

endmodule

module niosII_scfifo_a341 (
	clock,
	q,
	full_dff,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	empty_dff,
	all_bits_transmitted,
	wrreq,
	data,
	comb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
output 	full_dff;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
output 	empty_dff;
input 	all_bits_transmitted;
input 	wrreq;
input 	[7:0] data;
input 	comb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_a_dpfifo_tq31 dpfifo(
	.clock(clock),
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.full_dff1(full_dff),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.r_sync_rst(r_sync_rst),
	.empty_dff1(empty_dff),
	.all_bits_transmitted(all_bits_transmitted),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.comb(comb),
	.GND_port(GND_port));

endmodule

module niosII_a_dpfifo_tq31 (
	clock,
	q,
	full_dff1,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	empty_dff1,
	all_bits_transmitted,
	wreq,
	data,
	comb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
output 	full_dff1;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
output 	empty_dff1;
input 	all_bits_transmitted;
input 	wreq;
input 	[7:0] data;
input 	comb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \wr_ptr|counter_reg_bit[6]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[5]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[5]~q ;
wire \ram_read_address[5]~5_combout ;
wire \low_addressa[6]~q ;
wire \ram_read_address[6]~6_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \low_addressa[5]~5_combout ;
wire \low_addressa[6]~6_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_will_be_2~0_combout ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \usedw_will_be_2~1_combout ;
wire \usedw_is_2_dff~q ;
wire \usedw_will_be_1~4_combout ;
wire \usedw_will_be_0~0_combout ;
wire \usedw_will_be_0~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~0_combout ;


niosII_altsyncram_dqb1 FIFOram(
	.clock0(clock),
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[6]~q ,\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_b({\ram_read_address[6]~6_combout ,\ram_read_address[5]~5_combout ,\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }));

niosII_cntr_0ab wr_ptr(
	.clock(clock),
	.full_dff(full_dff1),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\wr_ptr|counter_reg_bit[6]~q ),
	.r_sync_rst(r_sync_rst),
	.all_bits_transmitted(all_bits_transmitted),
	.GND_port(GND_port));

niosII_cntr_ca7 usedw_counter(
	.clock(clock),
	.full_dff(full_dff1),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.r_sync_rst(r_sync_rst),
	.all_bits_transmitted(all_bits_transmitted),
	.updown(wreq),
	.comb(comb),
	.GND_port(GND_port));

niosII_cntr_v9b rd_ptr_msb(
	.clock(clock),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.r_sync_rst(r_sync_rst),
	.comb(comb),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(comb),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

dffeas \low_addressa[5] (
	.clk(clock),
	.d(\low_addressa[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[5]~q ),
	.prn(vcc));
defparam \low_addressa[5] .is_wysiwyg = "true";
defparam \low_addressa[5] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[5]~5_combout ),
	.cout());
defparam \ram_read_address[5]~5 .lut_mask = 16'hAACC;
defparam \ram_read_address[5]~5 .sum_lutc_input = "datac";

dffeas \low_addressa[6] (
	.clk(clock),
	.d(\low_addressa[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[6]~q ),
	.prn(vcc));
defparam \low_addressa[6] .is_wysiwyg = "true";
defparam \low_addressa[6] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[6]~6_combout ),
	.cout());
defparam \ram_read_address[6]~6 .lut_mask = 16'hAACC;
defparam \ram_read_address[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(comb),
	.datac(\rd_ptr_lsb~q ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'h8BFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(r_sync_rst),
	.datab(\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'h7777;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(r_sync_rst),
	.datab(comb),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEEEE;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hACFF;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hACFF;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hACFF;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hACFF;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[5]~5_combout ),
	.cout());
defparam \low_addressa[5]~5 .lut_mask = 16'hACFF;
defparam \low_addressa[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[6]~6_combout ),
	.cout());
defparam \low_addressa[6]~6 .lut_mask = 16'hACFF;
defparam \low_addressa[6]~6 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \_~0 (
	.dataa(counter_reg_bit_6),
	.datab(counter_reg_bit_5),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_3),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFFE;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(counter_reg_bit_1),
	.datab(wreq),
	.datac(counter_reg_bit_2),
	.datad(\_~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(counter_reg_bit_0),
	.datab(full_dff1),
	.datac(comb),
	.datad(\_~1_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFFEF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_2~0 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(comb),
	.cin(gnd),
	.combout(\usedw_will_be_2~0_combout ),
	.cout());
defparam \usedw_will_be_2~0 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_6),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hEFFF;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~4 (
	.dataa(\_~3_combout ),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_2),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hBFFF;
defparam \_~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~1 (
	.dataa(\usedw_will_be_2~0_combout ),
	.datab(comb),
	.datac(\_~4_combout ),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_2~1_combout ),
	.cout());
defparam \usedw_will_be_2~1 .lut_mask = 16'hFEFF;
defparam \usedw_will_be_2~1 .sum_lutc_input = "datac";

dffeas usedw_is_2_dff(
	.clk(clock),
	.d(\usedw_will_be_2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_2_dff~q ),
	.prn(vcc));
defparam usedw_is_2_dff.is_wysiwyg = "true";
defparam usedw_is_2_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~4 (
	.dataa(all_bits_transmitted),
	.datab(full_dff1),
	.datac(comb),
	.datad(\usedw_is_2_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~4_combout ),
	.cout());
defparam \usedw_will_be_1~4 .lut_mask = 16'hFFFD;
defparam \usedw_will_be_1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(comb),
	.cin(gnd),
	.combout(\usedw_will_be_0~0_combout ),
	.cout());
defparam \usedw_will_be_0~0 .lut_mask = 16'hBFEF;
defparam \usedw_will_be_0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~1 (
	.dataa(\usedw_will_be_0~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\usedw_will_be_0~1_combout ),
	.cout());
defparam \usedw_will_be_0~1 .lut_mask = 16'hAAFF;
defparam \usedw_will_be_0~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\usedw_will_be_0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(wreq),
	.datac(comb),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBEFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(\usedw_will_be_1~4_combout ),
	.datab(\usedw_will_be_1~2_combout ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hEEFF;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(r_sync_rst),
	.datab(wreq),
	.datac(\usedw_will_be_1~3_combout ),
	.datad(\usedw_will_be_0~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hFF7F;
defparam \empty_dff~0 .sum_lutc_input = "datac";

endmodule

module niosII_altsyncram_dqb1 (
	clock0,
	q_b,
	address_a,
	wren_a,
	data_a,
	address_b)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[7:0] q_b;
input 	[6:0] address_a;
input 	wren_a;
input 	[7:0] data_a;
input 	[6:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module niosII_cntr_0ab (
	clock,
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	r_sync_rst,
	all_bits_transmitted,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	r_sync_rst;
input 	all_bits_transmitted;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(r_sync_rst),
	.datab(all_bits_transmitted),
	.datac(gnd),
	.datad(full_dff),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hEEFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module niosII_cntr_ca7 (
	clock,
	full_dff,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	all_bits_transmitted,
	updown,
	comb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	full_dff;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
input 	all_bits_transmitted;
input 	updown;
input 	comb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;
wire \_~2_combout ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A6F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(all_bits_transmitted),
	.datab(full_dff),
	.datac(r_sync_rst),
	.datad(comb),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hF9F6;
defparam \_~2 .sum_lutc_input = "datac";

endmodule

module niosII_cntr_v9b (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	r_sync_rst,
	comb,
	rd_ptr_lsb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	r_sync_rst;
input 	comb;
input 	rd_ptr_lsb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(r_sync_rst),
	.datab(comb),
	.datac(gnd),
	.datad(rd_ptr_lsb),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hEEFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_altera_up_rs232_out_serializer (
	wire_pll7_clk_0,
	write_fifo_write_en,
	fifo_write_space_7,
	fifo_write_space_6,
	fifo_write_space_5,
	fifo_write_space_4,
	fifo_write_space_3,
	fifo_write_space_2,
	fifo_write_space_1,
	fifo_write_space_0,
	serial_data_out1,
	r_sync_rst,
	data_to_uart_0,
	data_to_uart_1,
	data_to_uart_2,
	data_to_uart_3,
	data_to_uart_4,
	data_to_uart_5,
	data_to_uart_6,
	data_to_uart_7,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	write_fifo_write_en;
output 	fifo_write_space_7;
output 	fifo_write_space_6;
output 	fifo_write_space_5;
output 	fifo_write_space_4;
output 	fifo_write_space_3;
output 	fifo_write_space_2;
output 	fifo_write_space_1;
output 	fifo_write_space_0;
output 	serial_data_out1;
input 	r_sync_rst;
input 	data_to_uart_0;
input 	data_to_uart_1;
input 	data_to_uart_2;
input 	data_to_uart_3;
input 	data_to_uart_4;
input 	data_to_uart_5;
input 	data_to_uart_6;
input 	data_to_uart_7;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \RS232_Out_Counters|baud_clock_rising_edge~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \RS232_Out_Counters|all_bits_transmitted~q ;
wire \comb~0_combout ;
wire \data_out_shift_reg[5]~4_combout ;
wire \fifo_write_space[0]~9 ;
wire \fifo_write_space[1]~11 ;
wire \fifo_write_space[2]~13 ;
wire \fifo_write_space[3]~15 ;
wire \fifo_write_space[4]~17 ;
wire \fifo_write_space[5]~19 ;
wire \fifo_write_space[6]~21 ;
wire \fifo_write_space[7]~22_combout ;
wire \fifo_write_space[6]~20_combout ;
wire \fifo_write_space[5]~18_combout ;
wire \fifo_write_space[4]~16_combout ;
wire \fifo_write_space[3]~14_combout ;
wire \fifo_write_space[2]~12_combout ;
wire \fifo_write_space[1]~10_combout ;
wire \fifo_write_space[0]~8_combout ;
wire \transmitting_data~0_combout ;
wire \transmitting_data~q ;
wire \read_fifo_en~0_combout ;
wire \data_out_shift_reg~10_combout ;
wire \data_out_shift_reg[8]~q ;
wire \data_out_shift_reg~9_combout ;
wire \data_out_shift_reg[5]~2_combout ;
wire \data_out_shift_reg[7]~q ;
wire \data_out_shift_reg~8_combout ;
wire \data_out_shift_reg[6]~q ;
wire \data_out_shift_reg~7_combout ;
wire \data_out_shift_reg[5]~q ;
wire \data_out_shift_reg~6_combout ;
wire \data_out_shift_reg[4]~q ;
wire \data_out_shift_reg~5_combout ;
wire \data_out_shift_reg[3]~q ;
wire \data_out_shift_reg~3_combout ;
wire \data_out_shift_reg[2]~q ;
wire \data_out_shift_reg~1_combout ;
wire \data_out_shift_reg[1]~q ;
wire \data_out_shift_reg~0_combout ;
wire \data_out_shift_reg[0]~q ;
wire \serial_data_out~0_combout ;


niosII_altera_up_sync_fifo_1 RS232_Out_FIFO(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.q_b_0(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.q_b_1(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.counter_reg_bit_1(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_5(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.counter_reg_bit_3(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_6(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.counter_reg_bit_2(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_4(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.q_b_2(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.r_sync_rst(r_sync_rst),
	.empty_dff(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.read_fifo_en(\read_fifo_en~0_combout ),
	.comb(\comb~0_combout ),
	.data_to_uart_0(data_to_uart_0),
	.data_out_shift_reg_5(\data_out_shift_reg[5]~4_combout ),
	.data_to_uart_1(data_to_uart_1),
	.data_to_uart_2(data_to_uart_2),
	.data_to_uart_3(data_to_uart_3),
	.data_to_uart_4(data_to_uart_4),
	.data_to_uart_5(data_to_uart_5),
	.data_to_uart_6(data_to_uart_6),
	.data_to_uart_7(data_to_uart_7),
	.GND_port(GND_port));

niosII_altera_up_rs232_counters_1 RS232_Out_Counters(
	.clk(wire_pll7_clk_0),
	.transmitting_data(\transmitting_data~q ),
	.r_sync_rst(r_sync_rst),
	.baud_clock_rising_edge1(\RS232_Out_Counters|baud_clock_rising_edge~q ),
	.all_bits_transmitted1(\RS232_Out_Counters|all_bits_transmitted~q ));

cycloneive_lcell_comb \comb~0 (
	.dataa(write_fifo_write_en),
	.datab(gnd),
	.datac(gnd),
	.datad(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hAAFF;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg[5]~4 (
	.dataa(r_sync_rst),
	.datab(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datac(\RS232_Out_Counters|all_bits_transmitted~q ),
	.datad(\transmitting_data~q ),
	.cin(gnd),
	.combout(\data_out_shift_reg[5]~4_combout ),
	.cout());
defparam \data_out_shift_reg[5]~4 .lut_mask = 16'hEFFF;
defparam \data_out_shift_reg[5]~4 .sum_lutc_input = "datac";

dffeas \fifo_write_space[7] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_7),
	.prn(vcc));
defparam \fifo_write_space[7] .is_wysiwyg = "true";
defparam \fifo_write_space[7] .power_up = "low";

dffeas \fifo_write_space[6] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_6),
	.prn(vcc));
defparam \fifo_write_space[6] .is_wysiwyg = "true";
defparam \fifo_write_space[6] .power_up = "low";

dffeas \fifo_write_space[5] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_5),
	.prn(vcc));
defparam \fifo_write_space[5] .is_wysiwyg = "true";
defparam \fifo_write_space[5] .power_up = "low";

dffeas \fifo_write_space[4] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_4),
	.prn(vcc));
defparam \fifo_write_space[4] .is_wysiwyg = "true";
defparam \fifo_write_space[4] .power_up = "low";

dffeas \fifo_write_space[3] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_3),
	.prn(vcc));
defparam \fifo_write_space[3] .is_wysiwyg = "true";
defparam \fifo_write_space[3] .power_up = "low";

dffeas \fifo_write_space[2] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_2),
	.prn(vcc));
defparam \fifo_write_space[2] .is_wysiwyg = "true";
defparam \fifo_write_space[2] .power_up = "low";

dffeas \fifo_write_space[1] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_1),
	.prn(vcc));
defparam \fifo_write_space[1] .is_wysiwyg = "true";
defparam \fifo_write_space[1] .power_up = "low";

dffeas \fifo_write_space[0] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_0),
	.prn(vcc));
defparam \fifo_write_space[0] .is_wysiwyg = "true";
defparam \fifo_write_space[0] .power_up = "low";

dffeas serial_data_out(
	.clk(wire_pll7_clk_0),
	.d(\serial_data_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(serial_data_out1),
	.prn(vcc));
defparam serial_data_out.is_wysiwyg = "true";
defparam serial_data_out.power_up = "low";

cycloneive_lcell_comb \fifo_write_space[0]~8 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\fifo_write_space[0]~8_combout ),
	.cout(\fifo_write_space[0]~9 ));
defparam \fifo_write_space[0]~8 .lut_mask = 16'hAA55;
defparam \fifo_write_space[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_write_space[1]~10 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[0]~9 ),
	.combout(\fifo_write_space[1]~10_combout ),
	.cout(\fifo_write_space[1]~11 ));
defparam \fifo_write_space[1]~10 .lut_mask = 16'h5AAF;
defparam \fifo_write_space[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[2]~12 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[1]~11 ),
	.combout(\fifo_write_space[2]~12_combout ),
	.cout(\fifo_write_space[2]~13 ));
defparam \fifo_write_space[2]~12 .lut_mask = 16'h5A5F;
defparam \fifo_write_space[2]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[3]~14 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[2]~13 ),
	.combout(\fifo_write_space[3]~14_combout ),
	.cout(\fifo_write_space[3]~15 ));
defparam \fifo_write_space[3]~14 .lut_mask = 16'h5AAF;
defparam \fifo_write_space[3]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[4]~16 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[3]~15 ),
	.combout(\fifo_write_space[4]~16_combout ),
	.cout(\fifo_write_space[4]~17 ));
defparam \fifo_write_space[4]~16 .lut_mask = 16'h5A5F;
defparam \fifo_write_space[4]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[5]~18 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[4]~17 ),
	.combout(\fifo_write_space[5]~18_combout ),
	.cout(\fifo_write_space[5]~19 ));
defparam \fifo_write_space[5]~18 .lut_mask = 16'h5AAF;
defparam \fifo_write_space[5]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[6]~20 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[5]~19 ),
	.combout(\fifo_write_space[6]~20_combout ),
	.cout(\fifo_write_space[6]~21 ));
defparam \fifo_write_space[6]~20 .lut_mask = 16'h5A5F;
defparam \fifo_write_space[6]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[7]~22 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fifo_write_space[6]~21 ),
	.combout(\fifo_write_space[7]~22_combout ),
	.cout());
defparam \fifo_write_space[7]~22 .lut_mask = 16'h5A5A;
defparam \fifo_write_space[7]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \transmitting_data~0 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datab(\transmitting_data~q ),
	.datac(gnd),
	.datad(\RS232_Out_Counters|all_bits_transmitted~q ),
	.cin(gnd),
	.combout(\transmitting_data~0_combout ),
	.cout());
defparam \transmitting_data~0 .lut_mask = 16'hEEFF;
defparam \transmitting_data~0 .sum_lutc_input = "datac";

dffeas transmitting_data(
	.clk(wire_pll7_clk_0),
	.d(\transmitting_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\transmitting_data~q ),
	.prn(vcc));
defparam transmitting_data.is_wysiwyg = "true";
defparam transmitting_data.power_up = "low";

cycloneive_lcell_comb \read_fifo_en~0 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datab(gnd),
	.datac(\RS232_Out_Counters|all_bits_transmitted~q ),
	.datad(\transmitting_data~q ),
	.cin(gnd),
	.combout(\read_fifo_en~0_combout ),
	.cout());
defparam \read_fifo_en~0 .lut_mask = 16'hAFFF;
defparam \read_fifo_en~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg~10 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(\RS232_Out_Counters|baud_clock_rising_edge~q ),
	.datac(\data_out_shift_reg[8]~q ),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~10_combout ),
	.cout());
defparam \data_out_shift_reg~10 .lut_mask = 16'hFAFC;
defparam \data_out_shift_reg~10 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[8] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(vcc),
	.q(\data_out_shift_reg[8]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[8] .is_wysiwyg = "true";
defparam \data_out_shift_reg[8] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~9 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(\data_out_shift_reg[8]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~9_combout ),
	.cout());
defparam \data_out_shift_reg~9 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg[5]~2 (
	.dataa(r_sync_rst),
	.datab(\RS232_Out_Counters|baud_clock_rising_edge~q ),
	.datac(\read_fifo_en~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_out_shift_reg[5]~2_combout ),
	.cout());
defparam \data_out_shift_reg[5]~2 .lut_mask = 16'hFEFE;
defparam \data_out_shift_reg[5]~2 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[7] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[5]~2_combout ),
	.q(\data_out_shift_reg[7]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[7] .is_wysiwyg = "true";
defparam \data_out_shift_reg[7] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~8 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(\data_out_shift_reg[7]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~8_combout ),
	.cout());
defparam \data_out_shift_reg~8 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~8 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[6] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[5]~2_combout ),
	.q(\data_out_shift_reg[6]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[6] .is_wysiwyg = "true";
defparam \data_out_shift_reg[6] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~7 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datab(\data_out_shift_reg[6]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~7_combout ),
	.cout());
defparam \data_out_shift_reg~7 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~7 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[5] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[5]~2_combout ),
	.q(\data_out_shift_reg[5]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[5] .is_wysiwyg = "true";
defparam \data_out_shift_reg[5] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~6 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datab(\data_out_shift_reg[5]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~6_combout ),
	.cout());
defparam \data_out_shift_reg~6 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~6 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[4] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[5]~2_combout ),
	.q(\data_out_shift_reg[4]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[4] .is_wysiwyg = "true";
defparam \data_out_shift_reg[4] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~5 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(\data_out_shift_reg[4]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~5_combout ),
	.cout());
defparam \data_out_shift_reg~5 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~5 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[3] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[5]~2_combout ),
	.q(\data_out_shift_reg[3]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[3] .is_wysiwyg = "true";
defparam \data_out_shift_reg[3] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~3 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(\data_out_shift_reg[3]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~3_combout ),
	.cout());
defparam \data_out_shift_reg~3 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~3 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[2] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[5]~2_combout ),
	.q(\data_out_shift_reg[2]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[2] .is_wysiwyg = "true";
defparam \data_out_shift_reg[2] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~1 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\data_out_shift_reg[2]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~1_combout ),
	.cout());
defparam \data_out_shift_reg~1 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~1 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[1] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[5]~2_combout ),
	.q(\data_out_shift_reg[1]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[1] .is_wysiwyg = "true";
defparam \data_out_shift_reg[1] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~0 (
	.dataa(\data_out_shift_reg[1]~q ),
	.datab(\data_out_shift_reg[0]~q ),
	.datac(\RS232_Out_Counters|baud_clock_rising_edge~q ),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~0_combout ),
	.cout());
defparam \data_out_shift_reg~0 .lut_mask = 16'hACFF;
defparam \data_out_shift_reg~0 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[0] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(vcc),
	.q(\data_out_shift_reg[0]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[0] .is_wysiwyg = "true";
defparam \data_out_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \serial_data_out~0 (
	.dataa(r_sync_rst),
	.datab(\data_out_shift_reg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\serial_data_out~0_combout ),
	.cout());
defparam \serial_data_out~0 .lut_mask = 16'hEEEE;
defparam \serial_data_out~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_rs232_counters_1 (
	clk,
	transmitting_data,
	r_sync_rst,
	baud_clock_rising_edge1,
	all_bits_transmitted1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	transmitting_data;
input 	r_sync_rst;
output 	baud_clock_rising_edge1;
output 	all_bits_transmitted1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \baud_counter[0]~10_combout ;
wire \baud_counter[0]~12_combout ;
wire \baud_counter[0]~q ;
wire \baud_counter[0]~11 ;
wire \baud_counter[1]~13_combout ;
wire \baud_counter[1]~q ;
wire \baud_counter[1]~14 ;
wire \baud_counter[2]~15_combout ;
wire \baud_counter[2]~q ;
wire \baud_counter[2]~16 ;
wire \baud_counter[3]~17_combout ;
wire \baud_counter[3]~q ;
wire \Equal0~0_combout ;
wire \baud_counter[3]~18 ;
wire \baud_counter[4]~19_combout ;
wire \baud_counter[4]~q ;
wire \baud_counter[4]~20 ;
wire \baud_counter[5]~21_combout ;
wire \baud_counter[5]~q ;
wire \baud_counter[5]~22 ;
wire \baud_counter[6]~23_combout ;
wire \baud_counter[6]~q ;
wire \baud_counter[6]~24 ;
wire \baud_counter[7]~25_combout ;
wire \baud_counter[7]~q ;
wire \Equal0~1_combout ;
wire \baud_counter[7]~26 ;
wire \baud_counter[8]~27_combout ;
wire \baud_counter[8]~q ;
wire \baud_counter[8]~28 ;
wire \baud_counter[9]~29_combout ;
wire \baud_counter[9]~q ;
wire \Equal0~2_combout ;
wire \baud_clock_rising_edge~0_combout ;
wire \bit_counter[2]~0_combout ;
wire \bit_counter[0]~2_combout ;
wire \bit_counter[0]~q ;
wire \bit_counter[1]~3_combout ;
wire \bit_counter[1]~q ;
wire \Add1~0_combout ;
wire \bit_counter[2]~1_combout ;
wire \bit_counter[2]~q ;
wire \Add1~1_combout ;
wire \bit_counter[3]~4_combout ;
wire \bit_counter[3]~q ;
wire \Equal2~0_combout ;
wire \all_bits_transmitted~0_combout ;


dffeas baud_clock_rising_edge(
	.clk(clk),
	.d(\baud_clock_rising_edge~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(baud_clock_rising_edge1),
	.prn(vcc));
defparam baud_clock_rising_edge.is_wysiwyg = "true";
defparam baud_clock_rising_edge.power_up = "low";

dffeas all_bits_transmitted(
	.clk(clk),
	.d(\all_bits_transmitted~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(all_bits_transmitted1),
	.prn(vcc));
defparam all_bits_transmitted.is_wysiwyg = "true";
defparam all_bits_transmitted.power_up = "low";

cycloneive_lcell_comb \baud_counter[0]~10 (
	.dataa(\baud_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\baud_counter[0]~10_combout ),
	.cout(\baud_counter[0]~11 ));
defparam \baud_counter[0]~10 .lut_mask = 16'h55AA;
defparam \baud_counter[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[0]~12 (
	.dataa(transmitting_data),
	.datab(\Equal0~2_combout ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\baud_counter[0]~12_combout ),
	.cout());
defparam \baud_counter[0]~12 .lut_mask = 16'hFF77;
defparam \baud_counter[0]~12 .sum_lutc_input = "datac";

dffeas \baud_counter[0] (
	.clk(clk),
	.d(\baud_counter[0]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[0]~q ),
	.prn(vcc));
defparam \baud_counter[0] .is_wysiwyg = "true";
defparam \baud_counter[0] .power_up = "low";

cycloneive_lcell_comb \baud_counter[1]~13 (
	.dataa(\baud_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[0]~11 ),
	.combout(\baud_counter[1]~13_combout ),
	.cout(\baud_counter[1]~14 ));
defparam \baud_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \baud_counter[1]~13 .sum_lutc_input = "cin";

dffeas \baud_counter[1] (
	.clk(clk),
	.d(\baud_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[1]~q ),
	.prn(vcc));
defparam \baud_counter[1] .is_wysiwyg = "true";
defparam \baud_counter[1] .power_up = "low";

cycloneive_lcell_comb \baud_counter[2]~15 (
	.dataa(\baud_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[1]~14 ),
	.combout(\baud_counter[2]~15_combout ),
	.cout(\baud_counter[2]~16 ));
defparam \baud_counter[2]~15 .lut_mask = 16'h5AAF;
defparam \baud_counter[2]~15 .sum_lutc_input = "cin";

dffeas \baud_counter[2] (
	.clk(clk),
	.d(\baud_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[2]~q ),
	.prn(vcc));
defparam \baud_counter[2] .is_wysiwyg = "true";
defparam \baud_counter[2] .power_up = "low";

cycloneive_lcell_comb \baud_counter[3]~17 (
	.dataa(\baud_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[2]~16 ),
	.combout(\baud_counter[3]~17_combout ),
	.cout(\baud_counter[3]~18 ));
defparam \baud_counter[3]~17 .lut_mask = 16'h5A5F;
defparam \baud_counter[3]~17 .sum_lutc_input = "cin";

dffeas \baud_counter[3] (
	.clk(clk),
	.d(\baud_counter[3]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[3]~q ),
	.prn(vcc));
defparam \baud_counter[3] .is_wysiwyg = "true";
defparam \baud_counter[3] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\baud_counter[0]~q ),
	.datab(\baud_counter[1]~q ),
	.datac(\baud_counter[3]~q ),
	.datad(\baud_counter[2]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFEFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[4]~19 (
	.dataa(\baud_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[3]~18 ),
	.combout(\baud_counter[4]~19_combout ),
	.cout(\baud_counter[4]~20 ));
defparam \baud_counter[4]~19 .lut_mask = 16'h5AAF;
defparam \baud_counter[4]~19 .sum_lutc_input = "cin";

dffeas \baud_counter[4] (
	.clk(clk),
	.d(\baud_counter[4]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[4]~q ),
	.prn(vcc));
defparam \baud_counter[4] .is_wysiwyg = "true";
defparam \baud_counter[4] .power_up = "low";

cycloneive_lcell_comb \baud_counter[5]~21 (
	.dataa(\baud_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[4]~20 ),
	.combout(\baud_counter[5]~21_combout ),
	.cout(\baud_counter[5]~22 ));
defparam \baud_counter[5]~21 .lut_mask = 16'h5A5F;
defparam \baud_counter[5]~21 .sum_lutc_input = "cin";

dffeas \baud_counter[5] (
	.clk(clk),
	.d(\baud_counter[5]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[5]~q ),
	.prn(vcc));
defparam \baud_counter[5] .is_wysiwyg = "true";
defparam \baud_counter[5] .power_up = "low";

cycloneive_lcell_comb \baud_counter[6]~23 (
	.dataa(\baud_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[5]~22 ),
	.combout(\baud_counter[6]~23_combout ),
	.cout(\baud_counter[6]~24 ));
defparam \baud_counter[6]~23 .lut_mask = 16'h5AAF;
defparam \baud_counter[6]~23 .sum_lutc_input = "cin";

dffeas \baud_counter[6] (
	.clk(clk),
	.d(\baud_counter[6]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[6]~q ),
	.prn(vcc));
defparam \baud_counter[6] .is_wysiwyg = "true";
defparam \baud_counter[6] .power_up = "low";

cycloneive_lcell_comb \baud_counter[7]~25 (
	.dataa(\baud_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[6]~24 ),
	.combout(\baud_counter[7]~25_combout ),
	.cout(\baud_counter[7]~26 ));
defparam \baud_counter[7]~25 .lut_mask = 16'h5A5F;
defparam \baud_counter[7]~25 .sum_lutc_input = "cin";

dffeas \baud_counter[7] (
	.clk(clk),
	.d(\baud_counter[7]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[7]~q ),
	.prn(vcc));
defparam \baud_counter[7] .is_wysiwyg = "true";
defparam \baud_counter[7] .power_up = "low";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\baud_counter[4]~q ),
	.datab(\baud_counter[7]~q ),
	.datac(\baud_counter[5]~q ),
	.datad(\baud_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[8]~27 (
	.dataa(\baud_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[7]~26 ),
	.combout(\baud_counter[8]~27_combout ),
	.cout(\baud_counter[8]~28 ));
defparam \baud_counter[8]~27 .lut_mask = 16'h5AAF;
defparam \baud_counter[8]~27 .sum_lutc_input = "cin";

dffeas \baud_counter[8] (
	.clk(clk),
	.d(\baud_counter[8]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[8]~q ),
	.prn(vcc));
defparam \baud_counter[8] .is_wysiwyg = "true";
defparam \baud_counter[8] .power_up = "low";

cycloneive_lcell_comb \baud_counter[9]~29 (
	.dataa(\baud_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\baud_counter[8]~28 ),
	.combout(\baud_counter[9]~29_combout ),
	.cout());
defparam \baud_counter[9]~29 .lut_mask = 16'h5A5A;
defparam \baud_counter[9]~29 .sum_lutc_input = "cin";

dffeas \baud_counter[9] (
	.clk(clk),
	.d(\baud_counter[9]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[0]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[9]~q ),
	.prn(vcc));
defparam \baud_counter[9] .is_wysiwyg = "true";
defparam \baud_counter[9] .power_up = "low";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\baud_counter[8]~q ),
	.datad(\baud_counter[9]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEFFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_clock_rising_edge~0 (
	.dataa(r_sync_rst),
	.datab(\Equal0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\baud_clock_rising_edge~0_combout ),
	.cout());
defparam \baud_clock_rising_edge~0 .lut_mask = 16'h7777;
defparam \baud_clock_rising_edge~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[2]~0 (
	.dataa(transmitting_data),
	.datab(\Equal2~0_combout ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\bit_counter[2]~0_combout ),
	.cout());
defparam \bit_counter[2]~0 .lut_mask = 16'hEEFF;
defparam \bit_counter[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[0]~2 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\Equal0~2_combout ),
	.datac(\bit_counter[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\bit_counter[0]~2_combout ),
	.cout());
defparam \bit_counter[0]~2 .lut_mask = 16'hBEBE;
defparam \bit_counter[0]~2 .sum_lutc_input = "datac";

dffeas \bit_counter[0] (
	.clk(clk),
	.d(\bit_counter[0]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[0]~q ),
	.prn(vcc));
defparam \bit_counter[0] .is_wysiwyg = "true";
defparam \bit_counter[0] .power_up = "low";

cycloneive_lcell_comb \bit_counter[1]~3 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[1]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\bit_counter[1]~3_combout ),
	.cout());
defparam \bit_counter[1]~3 .lut_mask = 16'hEBBE;
defparam \bit_counter[1]~3 .sum_lutc_input = "datac";

dffeas \bit_counter[1] (
	.clk(clk),
	.d(\bit_counter[1]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[1]~q ),
	.prn(vcc));
defparam \bit_counter[1] .is_wysiwyg = "true";
defparam \bit_counter[1] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(\bit_counter[2]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'hC33C;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[2]~1 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[2]~q ),
	.datac(\Add1~0_combout ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\bit_counter[2]~1_combout ),
	.cout());
defparam \bit_counter[2]~1 .lut_mask = 16'hFAFC;
defparam \bit_counter[2]~1 .sum_lutc_input = "datac";

dffeas \bit_counter[2] (
	.clk(clk),
	.d(\bit_counter[2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[2]~q ),
	.prn(vcc));
defparam \bit_counter[2] .is_wysiwyg = "true";
defparam \bit_counter[2] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(\bit_counter[3]~q ),
	.datab(\bit_counter[2]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[3]~4 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[3]~q ),
	.datac(\Add1~1_combout ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\bit_counter[3]~4_combout ),
	.cout());
defparam \bit_counter[3]~4 .lut_mask = 16'hFAFC;
defparam \bit_counter[3]~4 .sum_lutc_input = "datac";

dffeas \bit_counter[3] (
	.clk(clk),
	.d(\bit_counter[3]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[3]~q ),
	.prn(vcc));
defparam \bit_counter[3] .is_wysiwyg = "true";
defparam \bit_counter[3] .power_up = "low";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(\bit_counter[2]~q ),
	.datab(\bit_counter[0]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hEFFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \all_bits_transmitted~0 (
	.dataa(r_sync_rst),
	.datab(\Equal2~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\all_bits_transmitted~0_combout ),
	.cout());
defparam \all_bits_transmitted~0 .lut_mask = 16'h7777;
defparam \all_bits_transmitted~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_sync_fifo_1 (
	wire_pll7_clk_0,
	q_b_0,
	write_fifo_write_en,
	full_dff,
	q_b_1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_3,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_4,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	r_sync_rst,
	empty_dff,
	read_fifo_en,
	comb,
	data_to_uart_0,
	data_out_shift_reg_5,
	data_to_uart_1,
	data_to_uart_2,
	data_to_uart_3,
	data_to_uart_4,
	data_to_uart_5,
	data_to_uart_6,
	data_to_uart_7,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	q_b_0;
input 	write_fifo_write_en;
output 	full_dff;
output 	q_b_1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_3;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_4;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	r_sync_rst;
output 	empty_dff;
input 	read_fifo_en;
input 	comb;
input 	data_to_uart_0;
input 	data_out_shift_reg_5;
input 	data_to_uart_1;
input 	data_to_uart_2;
input 	data_to_uart_3;
input 	data_to_uart_4;
input 	data_to_uart_5;
input 	data_to_uart_6;
input 	data_to_uart_7;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_4 Sync_FIFO(
	.clock(wire_pll7_clk_0),
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(full_dff),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_4(counter_reg_bit_4),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.read_fifo_en(read_fifo_en),
	.wrreq(comb),
	.data({data_to_uart_7,data_to_uart_6,data_to_uart_5,data_to_uart_4,data_to_uart_3,data_to_uart_2,data_to_uart_1,data_to_uart_0}),
	.data_out_shift_reg_5(data_out_shift_reg_5),
	.GND_port(GND_port));

endmodule

module niosII_scfifo_4 (
	clock,
	q,
	write_fifo_write_en,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_3,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_4,
	r_sync_rst,
	empty_dff,
	read_fifo_en,
	wrreq,
	data,
	data_out_shift_reg_5,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
input 	write_fifo_write_en;
output 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_3;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_4;
input 	r_sync_rst;
output 	empty_dff;
input 	read_fifo_en;
input 	wrreq;
input 	[7:0] data;
input 	data_out_shift_reg_5;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_a341_1 auto_generated(
	.clock(clock),
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(full_dff),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_4(counter_reg_bit_4),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.read_fifo_en(read_fifo_en),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.data_out_shift_reg_5(data_out_shift_reg_5),
	.GND_port(GND_port));

endmodule

module niosII_scfifo_a341_1 (
	clock,
	q,
	write_fifo_write_en,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_3,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_4,
	r_sync_rst,
	empty_dff,
	read_fifo_en,
	wrreq,
	data,
	data_out_shift_reg_5,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
input 	write_fifo_write_en;
output 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_3;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_4;
input 	r_sync_rst;
output 	empty_dff;
input 	read_fifo_en;
input 	wrreq;
input 	[7:0] data;
input 	data_out_shift_reg_5;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_a_dpfifo_tq31_1 dpfifo(
	.clock(clock),
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff1(full_dff),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_4(counter_reg_bit_4),
	.r_sync_rst(r_sync_rst),
	.empty_dff1(empty_dff),
	.read_fifo_en(read_fifo_en),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.data_out_shift_reg_5(data_out_shift_reg_5),
	.GND_port(GND_port));

endmodule

module niosII_a_dpfifo_tq31_1 (
	clock,
	q,
	write_fifo_write_en,
	full_dff1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_3,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_4,
	r_sync_rst,
	empty_dff1,
	read_fifo_en,
	wreq,
	data,
	data_out_shift_reg_5,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
input 	write_fifo_write_en;
output 	full_dff1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_3;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_4;
input 	r_sync_rst;
output 	empty_dff1;
input 	read_fifo_en;
input 	wreq;
input 	[7:0] data;
input 	data_out_shift_reg_5;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \wr_ptr|counter_reg_bit[6]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[5]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[5]~q ;
wire \ram_read_address[5]~5_combout ;
wire \low_addressa[6]~q ;
wire \ram_read_address[6]~6_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \low_addressa[5]~5_combout ;
wire \low_addressa[6]~6_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_will_be_2~0_combout ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \usedw_will_be_2~1_combout ;
wire \usedw_is_2_dff~q ;
wire \usedw_will_be_1~4_combout ;
wire \usedw_will_be_0~0_combout ;
wire \usedw_will_be_0~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~0_combout ;


niosII_cntr_ca7_1 usedw_counter(
	.clock(clock),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(full_dff1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_4(counter_reg_bit_4),
	.r_sync_rst(r_sync_rst),
	.read_fifo_en(read_fifo_en),
	.updown(wreq),
	.GND_port(GND_port));

niosII_cntr_v9b_1 rd_ptr_msb(
	.clock(clock),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.r_sync_rst(r_sync_rst),
	.read_fifo_en(read_fifo_en),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port));

niosII_altsyncram_dqb1_1 FIFOram(
	.clock0(clock),
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[6]~q ,\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_b({\ram_read_address[6]~6_combout ,\ram_read_address[5]~5_combout ,\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }));

niosII_cntr_0ab_1 wr_ptr(
	.clock(clock),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(full_dff1),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\wr_ptr|counter_reg_bit[6]~q ),
	.r_sync_rst(r_sync_rst),
	.GND_port(GND_port));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_shift_reg_5),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(read_fifo_en),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

dffeas \low_addressa[5] (
	.clk(clock),
	.d(\low_addressa[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[5]~q ),
	.prn(vcc));
defparam \low_addressa[5] .is_wysiwyg = "true";
defparam \low_addressa[5] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[5]~5_combout ),
	.cout());
defparam \ram_read_address[5]~5 .lut_mask = 16'hAACC;
defparam \ram_read_address[5]~5 .sum_lutc_input = "datac";

dffeas \low_addressa[6] (
	.clk(clock),
	.d(\low_addressa[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[6]~q ),
	.prn(vcc));
defparam \low_addressa[6] .is_wysiwyg = "true";
defparam \low_addressa[6] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[6]~6_combout ),
	.cout());
defparam \ram_read_address[6]~6 .lut_mask = 16'hAACC;
defparam \ram_read_address[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(read_fifo_en),
	.datac(\rd_ptr_lsb~q ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'h8BFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(r_sync_rst),
	.datab(\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'h7777;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hACFF;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hACFF;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hACFF;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hACFF;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[5]~5_combout ),
	.cout());
defparam \low_addressa[5]~5 .lut_mask = 16'hACFF;
defparam \low_addressa[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[6]~6_combout ),
	.cout());
defparam \low_addressa[6]~6 .lut_mask = 16'hACFF;
defparam \low_addressa[6]~6 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \_~0 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_3),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFFE;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(write_fifo_write_en),
	.datab(counter_reg_bit_6),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(full_dff1),
	.datab(read_fifo_en),
	.datac(\_~0_combout ),
	.datad(\_~1_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFFFB;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_2~0 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\usedw_will_be_2~0_combout ),
	.cout());
defparam \usedw_will_be_2~0 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_6),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hEFFF;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~4 (
	.dataa(\_~3_combout ),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_3),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hBFFF;
defparam \_~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~1 (
	.dataa(\usedw_will_be_2~0_combout ),
	.datab(read_fifo_en),
	.datac(\_~4_combout ),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_2~1_combout ),
	.cout());
defparam \usedw_will_be_2~1 .lut_mask = 16'hFEFF;
defparam \usedw_will_be_2~1 .sum_lutc_input = "datac";

dffeas usedw_is_2_dff(
	.clk(clock),
	.d(\usedw_will_be_2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_2_dff~q ),
	.prn(vcc));
defparam usedw_is_2_dff.is_wysiwyg = "true";
defparam usedw_is_2_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~4 (
	.dataa(write_fifo_write_en),
	.datab(full_dff1),
	.datac(read_fifo_en),
	.datad(\usedw_is_2_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~4_combout ),
	.cout());
defparam \usedw_will_be_1~4 .lut_mask = 16'hFFFD;
defparam \usedw_will_be_1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\usedw_will_be_0~0_combout ),
	.cout());
defparam \usedw_will_be_0~0 .lut_mask = 16'hBFEF;
defparam \usedw_will_be_0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~1 (
	.dataa(\usedw_will_be_0~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\usedw_will_be_0~1_combout ),
	.cout());
defparam \usedw_will_be_0~1 .lut_mask = 16'hAAFF;
defparam \usedw_will_be_0~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\usedw_will_be_0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(wreq),
	.datac(read_fifo_en),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBEFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(\usedw_will_be_1~4_combout ),
	.datab(\usedw_will_be_1~2_combout ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hEEFF;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(r_sync_rst),
	.datab(wreq),
	.datac(\usedw_will_be_1~3_combout ),
	.datad(\usedw_will_be_0~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hFF7F;
defparam \empty_dff~0 .sum_lutc_input = "datac";

endmodule

module niosII_altsyncram_dqb1_1 (
	clock0,
	q_b,
	address_a,
	wren_a,
	data_a,
	address_b)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[7:0] q_b;
input 	[6:0] address_a;
input 	wren_a;
input 	[7:0] data_a;
input 	[6:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosII_rs232_0:rs232_0|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module niosII_cntr_0ab_1 (
	clock,
	write_fifo_write_en,
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	r_sync_rst,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	write_fifo_write_en;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	r_sync_rst;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(r_sync_rst),
	.datab(write_fifo_write_en),
	.datac(gnd),
	.datad(full_dff),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hEEFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module niosII_cntr_ca7_1 (
	clock,
	write_fifo_write_en,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_3,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_4,
	r_sync_rst,
	read_fifo_en,
	updown,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	write_fifo_write_en;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_3;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_4;
input 	r_sync_rst;
input 	read_fifo_en;
input 	updown;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(write_fifo_write_en),
	.datab(full_dff),
	.datac(r_sync_rst),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hF9F6;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A6F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module niosII_cntr_v9b_1 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	r_sync_rst,
	read_fifo_en,
	rd_ptr_lsb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	r_sync_rst;
input 	read_fifo_en;
input 	rd_ptr_lsb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(r_sync_rst),
	.datab(read_fifo_en),
	.datac(gnd),
	.datad(rd_ptr_lsb),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hEEFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_niosII_rs232_0_1 (
	wire_pll7_clk_0,
	W_alu_result_2,
	readdata_0,
	irq1,
	readdata_1,
	readdata_23,
	readdata_22,
	readdata_21,
	readdata_20,
	readdata_19,
	readdata_18,
	readdata_17,
	readdata_16,
	serial_data_out,
	r_sync_rst,
	cp_valid,
	data,
	data1,
	read_latency_shift_reg,
	data_to_uart_0,
	data2,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	data_to_uart_1,
	readdata_15,
	readdata_9,
	readdata_8,
	data_to_uart_2,
	comb,
	data_to_uart_3,
	data_to_uart_4,
	data_to_uart_5,
	data_to_uart_6,
	data_to_uart_7,
	GND_port,
	rs232_1_RXD)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_2;
output 	readdata_0;
output 	irq1;
output 	readdata_1;
output 	readdata_23;
output 	readdata_22;
output 	readdata_21;
output 	readdata_20;
output 	readdata_19;
output 	readdata_18;
output 	readdata_17;
output 	readdata_16;
output 	serial_data_out;
input 	r_sync_rst;
input 	cp_valid;
input 	data;
input 	data1;
input 	read_latency_shift_reg;
input 	data_to_uart_0;
input 	data2;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
input 	data_to_uart_1;
output 	readdata_15;
output 	readdata_9;
output 	readdata_8;
input 	data_to_uart_2;
input 	comb;
input 	data_to_uart_3;
input 	data_to_uart_4;
input 	data_to_uart_5;
input 	data_to_uart_6;
input 	data_to_uart_7;
input 	GND_port;
input 	rs232_1_RXD;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write_fifo_write_en~q ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \RS232_Out_Serializer|fifo_write_space[7]~q ;
wire \RS232_Out_Serializer|fifo_write_space[6]~q ;
wire \RS232_Out_Serializer|fifo_write_space[5]~q ;
wire \RS232_Out_Serializer|fifo_write_space[4]~q ;
wire \RS232_Out_Serializer|fifo_write_space[3]~q ;
wire \RS232_Out_Serializer|fifo_write_space[2]~q ;
wire \RS232_Out_Serializer|fifo_write_space[1]~q ;
wire \RS232_Out_Serializer|fifo_write_space[0]~q ;
wire \write_fifo_write_en~0_combout ;
wire \RS232_In_Deserializer|fifo_read_available[7]~q ;
wire \RS232_In_Deserializer|fifo_read_available[6]~q ;
wire \RS232_In_Deserializer|fifo_read_available[5]~q ;
wire \RS232_In_Deserializer|fifo_read_available[4]~q ;
wire \RS232_In_Deserializer|fifo_read_available[3]~q ;
wire \RS232_In_Deserializer|fifo_read_available[2]~q ;
wire \RS232_In_Deserializer|fifo_read_available[1]~q ;
wire \RS232_In_Deserializer|fifo_read_available[0]~q ;
wire \RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \write_interrupt_en~0_combout ;
wire \write_interrupt_en~1_combout ;
wire \read_interrupt_en~q ;
wire \readdata~0_combout ;
wire \readdata[19]~1_combout ;
wire \read_interrupt~0_combout ;
wire \read_interrupt~q ;
wire \write_interrupt_en~q ;
wire \write_interrupt~0_combout ;
wire \write_interrupt~q ;
wire \irq~0_combout ;
wire \readdata~2_combout ;
wire \readdata~9_combout ;
wire \readdata~10_combout ;
wire \readdata~11_combout ;
wire \readdata~12_combout ;
wire \readdata~13_combout ;
wire \readdata~14_combout ;
wire \readdata~15_combout ;
wire \readdata~16_combout ;
wire \readdata~3_combout ;
wire \readdata~4_combout ;
wire \readdata~5_combout ;
wire \readdata~6_combout ;
wire \readdata~7_combout ;
wire \readdata~8_combout ;
wire \readdata~17_combout ;
wire \readdata~18_combout ;
wire \readdata~19_combout ;


niosII_altera_up_rs232_in_deserializer_1 RS232_In_Deserializer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.W_alu_result_2(W_alu_result_2),
	.q_b_0(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.r_sync_rst(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.fifo_read_available_7(\RS232_In_Deserializer|fifo_read_available[7]~q ),
	.fifo_read_available_6(\RS232_In_Deserializer|fifo_read_available[6]~q ),
	.fifo_read_available_5(\RS232_In_Deserializer|fifo_read_available[5]~q ),
	.fifo_read_available_4(\RS232_In_Deserializer|fifo_read_available[4]~q ),
	.fifo_read_available_3(\RS232_In_Deserializer|fifo_read_available[3]~q ),
	.fifo_read_available_2(\RS232_In_Deserializer|fifo_read_available[2]~q ),
	.fifo_read_available_1(\RS232_In_Deserializer|fifo_read_available[1]~q ),
	.fifo_read_available_0(\RS232_In_Deserializer|fifo_read_available[0]~q ),
	.empty_dff(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.comb(comb),
	.GND_port(GND_port),
	.rs232_1_RXD(rs232_1_RXD));

niosII_altera_up_rs232_out_serializer_1 RS232_Out_Serializer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.write_fifo_write_en(\write_fifo_write_en~q ),
	.fifo_write_space_7(\RS232_Out_Serializer|fifo_write_space[7]~q ),
	.fifo_write_space_6(\RS232_Out_Serializer|fifo_write_space[6]~q ),
	.fifo_write_space_5(\RS232_Out_Serializer|fifo_write_space[5]~q ),
	.fifo_write_space_4(\RS232_Out_Serializer|fifo_write_space[4]~q ),
	.fifo_write_space_3(\RS232_Out_Serializer|fifo_write_space[3]~q ),
	.fifo_write_space_2(\RS232_Out_Serializer|fifo_write_space[2]~q ),
	.fifo_write_space_1(\RS232_Out_Serializer|fifo_write_space[1]~q ),
	.fifo_write_space_0(\RS232_Out_Serializer|fifo_write_space[0]~q ),
	.serial_data_out1(serial_data_out),
	.r_sync_rst(r_sync_rst),
	.data_to_uart_0(data_to_uart_0),
	.data_to_uart_1(data_to_uart_1),
	.data_to_uart_2(data_to_uart_2),
	.data_to_uart_3(data_to_uart_3),
	.data_to_uart_4(data_to_uart_4),
	.data_to_uart_5(data_to_uart_5),
	.data_to_uart_6(data_to_uart_6),
	.data_to_uart_7(data_to_uart_7),
	.GND_port(GND_port));

dffeas write_fifo_write_en(
	.clk(wire_pll7_clk_0),
	.d(\write_fifo_write_en~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\write_fifo_write_en~q ),
	.prn(vcc));
defparam write_fifo_write_en.is_wysiwyg = "true";
defparam write_fifo_write_en.power_up = "low";

cycloneive_lcell_comb \write_fifo_write_en~0 (
	.dataa(cp_valid),
	.datab(data2),
	.datac(read_latency_shift_reg),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\write_fifo_write_en~0_combout ),
	.cout());
defparam \write_fifo_write_en~0 .lut_mask = 16'hFEFF;
defparam \write_fifo_write_en~0 .sum_lutc_input = "datac";

dffeas \readdata[0] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas irq(
	.clk(wire_pll7_clk_0),
	.d(\irq~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(irq1),
	.prn(vcc));
defparam irq.is_wysiwyg = "true";
defparam irq.power_up = "low";

dffeas \readdata[1] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[23] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[22] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[21] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[20] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[19] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[18] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[17] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[16] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[2] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[15] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[9] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[8] (
	.clk(wire_pll7_clk_0),
	.d(\readdata~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[19]~1_combout ),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

cycloneive_lcell_comb \write_interrupt_en~0 (
	.dataa(cp_valid),
	.datab(W_alu_result_2),
	.datac(data2),
	.datad(read_latency_shift_reg),
	.cin(gnd),
	.combout(\write_interrupt_en~0_combout ),
	.cout());
defparam \write_interrupt_en~0 .lut_mask = 16'h7FFF;
defparam \write_interrupt_en~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_interrupt_en~1 (
	.dataa(\write_interrupt_en~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\write_interrupt_en~1_combout ),
	.cout());
defparam \write_interrupt_en~1 .lut_mask = 16'hFF55;
defparam \write_interrupt_en~1 .sum_lutc_input = "datac";

dffeas read_interrupt_en(
	.clk(wire_pll7_clk_0),
	.d(data),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_interrupt_en~1_combout ),
	.q(\read_interrupt_en~q ),
	.prn(vcc));
defparam read_interrupt_en.is_wysiwyg = "true";
defparam read_interrupt_en.power_up = "low";

cycloneive_lcell_comb \readdata~0 (
	.dataa(\read_interrupt_en~q ),
	.datab(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hAACC;
defparam \readdata~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[19]~1 (
	.dataa(gnd),
	.datab(cp_valid),
	.datac(read_latency_shift_reg),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata[19]~1_combout ),
	.cout());
defparam \readdata[19]~1 .lut_mask = 16'hFFFC;
defparam \readdata[19]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_interrupt~0 (
	.dataa(\read_interrupt_en~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[7]~q ),
	.datac(\RS232_In_Deserializer|fifo_read_available[6]~q ),
	.datad(\RS232_In_Deserializer|fifo_read_available[5]~q ),
	.cin(gnd),
	.combout(\read_interrupt~0_combout ),
	.cout());
defparam \read_interrupt~0 .lut_mask = 16'hFFFE;
defparam \read_interrupt~0 .sum_lutc_input = "datac";

dffeas read_interrupt(
	.clk(wire_pll7_clk_0),
	.d(\read_interrupt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\read_interrupt~q ),
	.prn(vcc));
defparam read_interrupt.is_wysiwyg = "true";
defparam read_interrupt.power_up = "low";

dffeas write_interrupt_en(
	.clk(wire_pll7_clk_0),
	.d(data1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_interrupt_en~1_combout ),
	.q(\write_interrupt_en~q ),
	.prn(vcc));
defparam write_interrupt_en.is_wysiwyg = "true";
defparam write_interrupt_en.power_up = "low";

cycloneive_lcell_comb \write_interrupt~0 (
	.dataa(\write_interrupt_en~q ),
	.datab(\RS232_Out_Serializer|fifo_write_space[7]~q ),
	.datac(\RS232_Out_Serializer|fifo_write_space[6]~q ),
	.datad(\RS232_Out_Serializer|fifo_write_space[5]~q ),
	.cin(gnd),
	.combout(\write_interrupt~0_combout ),
	.cout());
defparam \write_interrupt~0 .lut_mask = 16'hFFFE;
defparam \write_interrupt~0 .sum_lutc_input = "datac";

dffeas write_interrupt(
	.clk(wire_pll7_clk_0),
	.d(\write_interrupt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\write_interrupt~q ),
	.prn(vcc));
defparam write_interrupt.is_wysiwyg = "true";
defparam write_interrupt.power_up = "low";

cycloneive_lcell_comb \irq~0 (
	.dataa(\read_interrupt~q ),
	.datab(\write_interrupt~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\irq~0_combout ),
	.cout());
defparam \irq~0 .lut_mask = 16'hEEEE;
defparam \irq~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~2 (
	.dataa(\write_interrupt_en~q ),
	.datab(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hAACC;
defparam \readdata~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~9 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[7]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[7]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~9_combout ),
	.cout());
defparam \readdata~9 .lut_mask = 16'hAACC;
defparam \readdata~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~10 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[6]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[6]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~10_combout ),
	.cout());
defparam \readdata~10 .lut_mask = 16'hAACC;
defparam \readdata~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~11 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[5]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[5]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~11_combout ),
	.cout());
defparam \readdata~11 .lut_mask = 16'hAACC;
defparam \readdata~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~12 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[4]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[4]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~12_combout ),
	.cout());
defparam \readdata~12 .lut_mask = 16'hAACC;
defparam \readdata~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~13 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[3]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[3]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~13_combout ),
	.cout());
defparam \readdata~13 .lut_mask = 16'hAACC;
defparam \readdata~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~14 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[2]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[2]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~14_combout ),
	.cout());
defparam \readdata~14 .lut_mask = 16'hAACC;
defparam \readdata~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~15 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[1]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[1]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~15_combout ),
	.cout());
defparam \readdata~15 .lut_mask = 16'hAACC;
defparam \readdata~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~16 (
	.dataa(\RS232_Out_Serializer|fifo_write_space[0]~q ),
	.datab(\RS232_In_Deserializer|fifo_read_available[0]~q ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~16_combout ),
	.cout());
defparam \readdata~16 .lut_mask = 16'hAACC;
defparam \readdata~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~3 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hAFFF;
defparam \readdata~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~4 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hAFFF;
defparam \readdata~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~5 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hAFFF;
defparam \readdata~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~6 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hAFFF;
defparam \readdata~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~7 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hAFFF;
defparam \readdata~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~8 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hAFFF;
defparam \readdata~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~17 (
	.dataa(\RS232_In_Deserializer|RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datab(gnd),
	.datac(r_sync_rst),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\readdata~17_combout ),
	.cout());
defparam \readdata~17 .lut_mask = 16'hAFFF;
defparam \readdata~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~18 (
	.dataa(W_alu_result_2),
	.datab(\write_interrupt~q ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata~18_combout ),
	.cout());
defparam \readdata~18 .lut_mask = 16'hEEFF;
defparam \readdata~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~19 (
	.dataa(W_alu_result_2),
	.datab(\read_interrupt~q ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata~19_combout ),
	.cout());
defparam \readdata~19 .lut_mask = 16'hEEFF;
defparam \readdata~19 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_rs232_in_deserializer_1 (
	wire_pll7_clk_0,
	W_alu_result_2,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	r_sync_rst,
	read_latency_shift_reg,
	fifo_read_available_7,
	fifo_read_available_6,
	fifo_read_available_5,
	fifo_read_available_4,
	fifo_read_available_3,
	fifo_read_available_2,
	fifo_read_available_1,
	fifo_read_available_0,
	empty_dff,
	comb,
	GND_port,
	rs232_1_RXD)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_2;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	r_sync_rst;
input 	read_latency_shift_reg;
output 	fifo_read_available_7;
output 	fifo_read_available_6;
output 	fifo_read_available_5;
output 	fifo_read_available_4;
output 	fifo_read_available_3;
output 	fifo_read_available_2;
output 	fifo_read_available_1;
output 	fifo_read_available_0;
output 	empty_dff;
input 	comb;
input 	GND_port;
input 	rs232_1_RXD;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \RS232_In_Counters|baud_clock_falling_edge~q ;
wire \receiving_data~q ;
wire \RS232_In_Counters|all_bits_transmitted~q ;
wire \comb~0_combout ;
wire \data_in_shift_reg[1]~q ;
wire \comb~1_combout ;
wire \data_in_shift_reg[2]~q ;
wire \data_in_shift_reg[3]~q ;
wire \data_in_shift_reg[4]~q ;
wire \data_in_shift_reg[5]~q ;
wire \data_in_shift_reg[6]~q ;
wire \data_in_shift_reg[7]~q ;
wire \data_in_shift_reg[8]~q ;
wire \data_in_shift_reg~0_combout ;
wire \data_in_shift_reg[1]~1_combout ;
wire \data_in_shift_reg~2_combout ;
wire \data_in_shift_reg~3_combout ;
wire \data_in_shift_reg~4_combout ;
wire \data_in_shift_reg~5_combout ;
wire \data_in_shift_reg~6_combout ;
wire \data_in_shift_reg~7_combout ;
wire \data_in_shift_reg[9]~q ;
wire \data_in_shift_reg~8_combout ;
wire \data_in_shift_reg~9_combout ;
wire \receiving_data~0_combout ;
wire \fifo_read_available~0_combout ;
wire \fifo_read_available~1_combout ;
wire \fifo_read_available~2_combout ;
wire \fifo_read_available~3_combout ;
wire \fifo_read_available~4_combout ;
wire \fifo_read_available~5_combout ;
wire \fifo_read_available~6_combout ;
wire \fifo_read_available~7_combout ;


niosII_altera_up_sync_fifo_2 RS232_In_FIFO(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.full_dff(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.counter_reg_bit_6(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.counter_reg_bit_5(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.all_bits_transmitted(\RS232_In_Counters|all_bits_transmitted~q ),
	.comb(\comb~0_combout ),
	.data_in_shift_reg_1(\data_in_shift_reg[1]~q ),
	.comb1(\comb~1_combout ),
	.data_in_shift_reg_2(\data_in_shift_reg[2]~q ),
	.data_in_shift_reg_3(\data_in_shift_reg[3]~q ),
	.data_in_shift_reg_4(\data_in_shift_reg[4]~q ),
	.data_in_shift_reg_5(\data_in_shift_reg[5]~q ),
	.data_in_shift_reg_6(\data_in_shift_reg[6]~q ),
	.data_in_shift_reg_7(\data_in_shift_reg[7]~q ),
	.data_in_shift_reg_8(\data_in_shift_reg[8]~q ),
	.GND_port(GND_port));

niosII_altera_up_rs232_counters_2 RS232_In_Counters(
	.clk(wire_pll7_clk_0),
	.baud_clock_falling_edge1(\RS232_In_Counters|baud_clock_falling_edge~q ),
	.receiving_data(\receiving_data~q ),
	.r_sync_rst(r_sync_rst),
	.all_bits_transmitted1(\RS232_In_Counters|all_bits_transmitted~q ));

dffeas receiving_data(
	.clk(wire_pll7_clk_0),
	.d(\receiving_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\receiving_data~q ),
	.prn(vcc));
defparam receiving_data.is_wysiwyg = "true";
defparam receiving_data.power_up = "low";

cycloneive_lcell_comb \comb~0 (
	.dataa(\RS232_In_Counters|all_bits_transmitted~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hAAFF;
defparam \comb~0 .sum_lutc_input = "datac";

dffeas \data_in_shift_reg[1] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[1]~1_combout ),
	.q(\data_in_shift_reg[1]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[1] .is_wysiwyg = "true";
defparam \data_in_shift_reg[1] .power_up = "low";

cycloneive_lcell_comb \comb~1 (
	.dataa(read_latency_shift_reg),
	.datab(empty_dff),
	.datac(comb),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\comb~1_combout ),
	.cout());
defparam \comb~1 .lut_mask = 16'hFEFF;
defparam \comb~1 .sum_lutc_input = "datac";

dffeas \data_in_shift_reg[2] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[1]~1_combout ),
	.q(\data_in_shift_reg[2]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[2] .is_wysiwyg = "true";
defparam \data_in_shift_reg[2] .power_up = "low";

dffeas \data_in_shift_reg[3] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[1]~1_combout ),
	.q(\data_in_shift_reg[3]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[3] .is_wysiwyg = "true";
defparam \data_in_shift_reg[3] .power_up = "low";

dffeas \data_in_shift_reg[4] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[1]~1_combout ),
	.q(\data_in_shift_reg[4]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[4] .is_wysiwyg = "true";
defparam \data_in_shift_reg[4] .power_up = "low";

dffeas \data_in_shift_reg[5] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[1]~1_combout ),
	.q(\data_in_shift_reg[5]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[5] .is_wysiwyg = "true";
defparam \data_in_shift_reg[5] .power_up = "low";

dffeas \data_in_shift_reg[6] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[1]~1_combout ),
	.q(\data_in_shift_reg[6]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[6] .is_wysiwyg = "true";
defparam \data_in_shift_reg[6] .power_up = "low";

dffeas \data_in_shift_reg[7] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[1]~1_combout ),
	.q(\data_in_shift_reg[7]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[7] .is_wysiwyg = "true";
defparam \data_in_shift_reg[7] .power_up = "low";

dffeas \data_in_shift_reg[8] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[1]~1_combout ),
	.q(\data_in_shift_reg[8]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[8] .is_wysiwyg = "true";
defparam \data_in_shift_reg[8] .power_up = "low";

cycloneive_lcell_comb \data_in_shift_reg~0 (
	.dataa(\data_in_shift_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~0_combout ),
	.cout());
defparam \data_in_shift_reg~0 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg[1]~1 (
	.dataa(r_sync_rst),
	.datab(\RS232_In_Counters|baud_clock_falling_edge~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_shift_reg[1]~1_combout ),
	.cout());
defparam \data_in_shift_reg[1]~1 .lut_mask = 16'hEEEE;
defparam \data_in_shift_reg[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~2 (
	.dataa(\data_in_shift_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~2_combout ),
	.cout());
defparam \data_in_shift_reg~2 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~3 (
	.dataa(\data_in_shift_reg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~3_combout ),
	.cout());
defparam \data_in_shift_reg~3 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~4 (
	.dataa(\data_in_shift_reg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~4_combout ),
	.cout());
defparam \data_in_shift_reg~4 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~5 (
	.dataa(\data_in_shift_reg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~5_combout ),
	.cout());
defparam \data_in_shift_reg~5 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~6 (
	.dataa(\data_in_shift_reg[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~6_combout ),
	.cout());
defparam \data_in_shift_reg~6 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~7 (
	.dataa(\data_in_shift_reg[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~7_combout ),
	.cout());
defparam \data_in_shift_reg~7 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~7 .sum_lutc_input = "datac";

dffeas \data_in_shift_reg[9] (
	.clk(wire_pll7_clk_0),
	.d(\data_in_shift_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[1]~1_combout ),
	.q(\data_in_shift_reg[9]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[9] .is_wysiwyg = "true";
defparam \data_in_shift_reg[9] .power_up = "low";

cycloneive_lcell_comb \data_in_shift_reg~8 (
	.dataa(\data_in_shift_reg[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~8_combout ),
	.cout());
defparam \data_in_shift_reg~8 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~9 (
	.dataa(rs232_1_RXD),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\data_in_shift_reg~9_combout ),
	.cout());
defparam \data_in_shift_reg~9 .lut_mask = 16'hAAFF;
defparam \data_in_shift_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \receiving_data~0 (
	.dataa(\receiving_data~q ),
	.datab(gnd),
	.datac(rs232_1_RXD),
	.datad(\RS232_In_Counters|all_bits_transmitted~q ),
	.cin(gnd),
	.combout(\receiving_data~0_combout ),
	.cout());
defparam \receiving_data~0 .lut_mask = 16'hAFFF;
defparam \receiving_data~0 .sum_lutc_input = "datac";

dffeas \fifo_read_available[7] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_7),
	.prn(vcc));
defparam \fifo_read_available[7] .is_wysiwyg = "true";
defparam \fifo_read_available[7] .power_up = "low";

dffeas \fifo_read_available[6] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_6),
	.prn(vcc));
defparam \fifo_read_available[6] .is_wysiwyg = "true";
defparam \fifo_read_available[6] .power_up = "low";

dffeas \fifo_read_available[5] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_5),
	.prn(vcc));
defparam \fifo_read_available[5] .is_wysiwyg = "true";
defparam \fifo_read_available[5] .power_up = "low";

dffeas \fifo_read_available[4] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_4),
	.prn(vcc));
defparam \fifo_read_available[4] .is_wysiwyg = "true";
defparam \fifo_read_available[4] .power_up = "low";

dffeas \fifo_read_available[3] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_3),
	.prn(vcc));
defparam \fifo_read_available[3] .is_wysiwyg = "true";
defparam \fifo_read_available[3] .power_up = "low";

dffeas \fifo_read_available[2] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_2),
	.prn(vcc));
defparam \fifo_read_available[2] .is_wysiwyg = "true";
defparam \fifo_read_available[2] .power_up = "low";

dffeas \fifo_read_available[1] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_1),
	.prn(vcc));
defparam \fifo_read_available[1] .is_wysiwyg = "true";
defparam \fifo_read_available[1] .power_up = "low";

dffeas \fifo_read_available[0] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_read_available~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_read_available_0),
	.prn(vcc));
defparam \fifo_read_available[0] .is_wysiwyg = "true";
defparam \fifo_read_available[0] .power_up = "low";

cycloneive_lcell_comb \fifo_read_available~0 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~0_combout ),
	.cout());
defparam \fifo_read_available~0 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~1 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~1_combout ),
	.cout());
defparam \fifo_read_available~1 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~2 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~2_combout ),
	.cout());
defparam \fifo_read_available~2 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~3 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~3_combout ),
	.cout());
defparam \fifo_read_available~3 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~4 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~4_combout ),
	.cout());
defparam \fifo_read_available~4 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~5 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~5_combout ),
	.cout());
defparam \fifo_read_available~5 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~6 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~6_combout ),
	.cout());
defparam \fifo_read_available~6 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_read_available~7 (
	.dataa(\RS232_In_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\fifo_read_available~7_combout ),
	.cout());
defparam \fifo_read_available~7 .lut_mask = 16'hAAFF;
defparam \fifo_read_available~7 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_rs232_counters_2 (
	clk,
	baud_clock_falling_edge1,
	receiving_data,
	r_sync_rst,
	all_bits_transmitted1)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	baud_clock_falling_edge1;
input 	receiving_data;
input 	r_sync_rst;
output 	all_bits_transmitted1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \baud_counter[0]~10_combout ;
wire \baud_counter[5]~22 ;
wire \baud_counter[6]~23_combout ;
wire \baud_counter[6]~q ;
wire \Equal0~0_combout ;
wire \baud_counter[6]~24 ;
wire \baud_counter[7]~25_combout ;
wire \baud_counter[7]~q ;
wire \baud_counter[7]~26 ;
wire \baud_counter[8]~27_combout ;
wire \baud_counter[8]~q ;
wire \baud_counter[8]~28 ;
wire \baud_counter[9]~29_combout ;
wire \baud_counter[9]~q ;
wire \Equal0~1_combout ;
wire \baud_counter[5]~14_combout ;
wire \baud_counter[0]~q ;
wire \baud_counter[0]~11 ;
wire \baud_counter[1]~12_combout ;
wire \baud_counter[1]~q ;
wire \baud_counter[1]~13 ;
wire \baud_counter[2]~15_combout ;
wire \baud_counter[2]~q ;
wire \baud_counter[2]~16 ;
wire \baud_counter[3]~17_combout ;
wire \baud_counter[3]~q ;
wire \baud_counter[3]~18 ;
wire \baud_counter[4]~19_combout ;
wire \baud_counter[4]~q ;
wire \baud_counter[4]~20 ;
wire \baud_counter[5]~21_combout ;
wire \baud_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \Equal1~2_combout ;
wire \bit_counter[2]~0_combout ;
wire \bit_counter[0]~2_combout ;
wire \bit_counter[0]~q ;
wire \bit_counter[1]~3_combout ;
wire \bit_counter[1]~q ;
wire \Add1~0_combout ;
wire \bit_counter[2]~1_combout ;
wire \bit_counter[2]~q ;
wire \Add1~1_combout ;
wire \bit_counter[3]~4_combout ;
wire \bit_counter[3]~q ;
wire \Equal2~0_combout ;
wire \all_bits_transmitted~0_combout ;


dffeas baud_clock_falling_edge(
	.clk(clk),
	.d(\Equal1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(baud_clock_falling_edge1),
	.prn(vcc));
defparam baud_clock_falling_edge.is_wysiwyg = "true";
defparam baud_clock_falling_edge.power_up = "low";

dffeas all_bits_transmitted(
	.clk(clk),
	.d(\all_bits_transmitted~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(all_bits_transmitted1),
	.prn(vcc));
defparam all_bits_transmitted.is_wysiwyg = "true";
defparam all_bits_transmitted.power_up = "low";

cycloneive_lcell_comb \baud_counter[0]~10 (
	.dataa(\baud_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\baud_counter[0]~10_combout ),
	.cout(\baud_counter[0]~11 ));
defparam \baud_counter[0]~10 .lut_mask = 16'h55AA;
defparam \baud_counter[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[5]~21 (
	.dataa(\baud_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[4]~20 ),
	.combout(\baud_counter[5]~21_combout ),
	.cout(\baud_counter[5]~22 ));
defparam \baud_counter[5]~21 .lut_mask = 16'h5A5F;
defparam \baud_counter[5]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \baud_counter[6]~23 (
	.dataa(\baud_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[5]~22 ),
	.combout(\baud_counter[6]~23_combout ),
	.cout(\baud_counter[6]~24 ));
defparam \baud_counter[6]~23 .lut_mask = 16'h5AAF;
defparam \baud_counter[6]~23 .sum_lutc_input = "cin";

dffeas \baud_counter[6] (
	.clk(clk),
	.d(\baud_counter[6]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[6]~q ),
	.prn(vcc));
defparam \baud_counter[6] .is_wysiwyg = "true";
defparam \baud_counter[6] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\baud_counter[1]~q ),
	.datab(\baud_counter[4]~q ),
	.datac(\baud_counter[2]~q ),
	.datad(\baud_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[7]~25 (
	.dataa(\baud_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[6]~24 ),
	.combout(\baud_counter[7]~25_combout ),
	.cout(\baud_counter[7]~26 ));
defparam \baud_counter[7]~25 .lut_mask = 16'h5A5F;
defparam \baud_counter[7]~25 .sum_lutc_input = "cin";

dffeas \baud_counter[7] (
	.clk(clk),
	.d(\baud_counter[7]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[7]~q ),
	.prn(vcc));
defparam \baud_counter[7] .is_wysiwyg = "true";
defparam \baud_counter[7] .power_up = "low";

cycloneive_lcell_comb \baud_counter[8]~27 (
	.dataa(\baud_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[7]~26 ),
	.combout(\baud_counter[8]~27_combout ),
	.cout(\baud_counter[8]~28 ));
defparam \baud_counter[8]~27 .lut_mask = 16'h5AAF;
defparam \baud_counter[8]~27 .sum_lutc_input = "cin";

dffeas \baud_counter[8] (
	.clk(clk),
	.d(\baud_counter[8]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[8]~q ),
	.prn(vcc));
defparam \baud_counter[8] .is_wysiwyg = "true";
defparam \baud_counter[8] .power_up = "low";

cycloneive_lcell_comb \baud_counter[9]~29 (
	.dataa(\baud_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\baud_counter[8]~28 ),
	.combout(\baud_counter[9]~29_combout ),
	.cout());
defparam \baud_counter[9]~29 .lut_mask = 16'h5A5A;
defparam \baud_counter[9]~29 .sum_lutc_input = "cin";

dffeas \baud_counter[9] (
	.clk(clk),
	.d(\baud_counter[9]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[9]~q ),
	.prn(vcc));
defparam \baud_counter[9] .is_wysiwyg = "true";
defparam \baud_counter[9] .power_up = "low";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\Equal0~0_combout ),
	.datab(\baud_counter[7]~q ),
	.datac(\Equal1~0_combout ),
	.datad(\baud_counter[9]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[5]~14 (
	.dataa(\Equal0~1_combout ),
	.datab(receiving_data),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\baud_counter[5]~14_combout ),
	.cout());
defparam \baud_counter[5]~14 .lut_mask = 16'hFF77;
defparam \baud_counter[5]~14 .sum_lutc_input = "datac";

dffeas \baud_counter[0] (
	.clk(clk),
	.d(\baud_counter[0]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[0]~q ),
	.prn(vcc));
defparam \baud_counter[0] .is_wysiwyg = "true";
defparam \baud_counter[0] .power_up = "low";

cycloneive_lcell_comb \baud_counter[1]~12 (
	.dataa(\baud_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[0]~11 ),
	.combout(\baud_counter[1]~12_combout ),
	.cout(\baud_counter[1]~13 ));
defparam \baud_counter[1]~12 .lut_mask = 16'h5A5F;
defparam \baud_counter[1]~12 .sum_lutc_input = "cin";

dffeas \baud_counter[1] (
	.clk(clk),
	.d(\baud_counter[1]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[1]~q ),
	.prn(vcc));
defparam \baud_counter[1] .is_wysiwyg = "true";
defparam \baud_counter[1] .power_up = "low";

cycloneive_lcell_comb \baud_counter[2]~15 (
	.dataa(\baud_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[1]~13 ),
	.combout(\baud_counter[2]~15_combout ),
	.cout(\baud_counter[2]~16 ));
defparam \baud_counter[2]~15 .lut_mask = 16'h5AAF;
defparam \baud_counter[2]~15 .sum_lutc_input = "cin";

dffeas \baud_counter[2] (
	.clk(clk),
	.d(\baud_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[2]~q ),
	.prn(vcc));
defparam \baud_counter[2] .is_wysiwyg = "true";
defparam \baud_counter[2] .power_up = "low";

cycloneive_lcell_comb \baud_counter[3]~17 (
	.dataa(\baud_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[2]~16 ),
	.combout(\baud_counter[3]~17_combout ),
	.cout(\baud_counter[3]~18 ));
defparam \baud_counter[3]~17 .lut_mask = 16'h5A5F;
defparam \baud_counter[3]~17 .sum_lutc_input = "cin";

dffeas \baud_counter[3] (
	.clk(clk),
	.d(\baud_counter[3]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[3]~q ),
	.prn(vcc));
defparam \baud_counter[3] .is_wysiwyg = "true";
defparam \baud_counter[3] .power_up = "low";

cycloneive_lcell_comb \baud_counter[4]~19 (
	.dataa(\baud_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[3]~18 ),
	.combout(\baud_counter[4]~19_combout ),
	.cout(\baud_counter[4]~20 ));
defparam \baud_counter[4]~19 .lut_mask = 16'h5AAF;
defparam \baud_counter[4]~19 .sum_lutc_input = "cin";

dffeas \baud_counter[4] (
	.clk(clk),
	.d(\baud_counter[4]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[4]~q ),
	.prn(vcc));
defparam \baud_counter[4] .is_wysiwyg = "true";
defparam \baud_counter[4] .power_up = "low";

dffeas \baud_counter[5] (
	.clk(clk),
	.d(\baud_counter[5]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[5]~14_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[5]~q ),
	.prn(vcc));
defparam \baud_counter[5] .is_wysiwyg = "true";
defparam \baud_counter[5] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\baud_counter[5]~q ),
	.datab(\baud_counter[8]~q ),
	.datac(\baud_counter[0]~q ),
	.datad(\baud_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(\baud_counter[1]~q ),
	.datab(\baud_counter[4]~q ),
	.datac(\baud_counter[2]~q ),
	.datad(\baud_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hEFFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(\Equal1~0_combout ),
	.datab(\baud_counter[7]~q ),
	.datac(\Equal1~1_combout ),
	.datad(\baud_counter[9]~q ),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'hFEFF;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[2]~0 (
	.dataa(\Equal2~0_combout ),
	.datab(receiving_data),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\bit_counter[2]~0_combout ),
	.cout());
defparam \bit_counter[2]~0 .lut_mask = 16'hEEFF;
defparam \bit_counter[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[0]~2 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[0]~q ),
	.datac(\Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\bit_counter[0]~2_combout ),
	.cout());
defparam \bit_counter[0]~2 .lut_mask = 16'hBEBE;
defparam \bit_counter[0]~2 .sum_lutc_input = "datac";

dffeas \bit_counter[0] (
	.clk(clk),
	.d(\bit_counter[0]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[0]~q ),
	.prn(vcc));
defparam \bit_counter[0] .is_wysiwyg = "true";
defparam \bit_counter[0] .power_up = "low";

cycloneive_lcell_comb \bit_counter[1]~3 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[1]~q ),
	.datac(\Equal0~1_combout ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\bit_counter[1]~3_combout ),
	.cout());
defparam \bit_counter[1]~3 .lut_mask = 16'hEBBE;
defparam \bit_counter[1]~3 .sum_lutc_input = "datac";

dffeas \bit_counter[1] (
	.clk(clk),
	.d(\bit_counter[1]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[1]~q ),
	.prn(vcc));
defparam \bit_counter[1] .is_wysiwyg = "true";
defparam \bit_counter[1] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(\bit_counter[2]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'hC33C;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[2]~1 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[2]~q ),
	.datac(\Add1~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\bit_counter[2]~1_combout ),
	.cout());
defparam \bit_counter[2]~1 .lut_mask = 16'hFAFC;
defparam \bit_counter[2]~1 .sum_lutc_input = "datac";

dffeas \bit_counter[2] (
	.clk(clk),
	.d(\bit_counter[2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[2]~q ),
	.prn(vcc));
defparam \bit_counter[2] .is_wysiwyg = "true";
defparam \bit_counter[2] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(\bit_counter[3]~q ),
	.datab(\bit_counter[2]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[3]~4 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[3]~q ),
	.datac(\Add1~1_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\bit_counter[3]~4_combout ),
	.cout());
defparam \bit_counter[3]~4 .lut_mask = 16'hFAFC;
defparam \bit_counter[3]~4 .sum_lutc_input = "datac";

dffeas \bit_counter[3] (
	.clk(clk),
	.d(\bit_counter[3]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[3]~q ),
	.prn(vcc));
defparam \bit_counter[3] .is_wysiwyg = "true";
defparam \bit_counter[3] .power_up = "low";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(\bit_counter[2]~q ),
	.datab(\bit_counter[0]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hEFFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \all_bits_transmitted~0 (
	.dataa(r_sync_rst),
	.datab(\Equal2~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\all_bits_transmitted~0_combout ),
	.cout());
defparam \all_bits_transmitted~0 .lut_mask = 16'h7777;
defparam \all_bits_transmitted~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_sync_fifo_2 (
	wire_pll7_clk_0,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	full_dff,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	empty_dff,
	all_bits_transmitted,
	comb,
	data_in_shift_reg_1,
	comb1,
	data_in_shift_reg_2,
	data_in_shift_reg_3,
	data_in_shift_reg_4,
	data_in_shift_reg_5,
	data_in_shift_reg_6,
	data_in_shift_reg_7,
	data_in_shift_reg_8,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	full_dff;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
output 	empty_dff;
input 	all_bits_transmitted;
input 	comb;
input 	data_in_shift_reg_1;
input 	comb1;
input 	data_in_shift_reg_2;
input 	data_in_shift_reg_3;
input 	data_in_shift_reg_4;
input 	data_in_shift_reg_5;
input 	data_in_shift_reg_6;
input 	data_in_shift_reg_7;
input 	data_in_shift_reg_8;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_5 Sync_FIFO(
	.clock(wire_pll7_clk_0),
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.full_dff(full_dff),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.all_bits_transmitted(all_bits_transmitted),
	.wrreq(comb),
	.data({data_in_shift_reg_8,data_in_shift_reg_7,data_in_shift_reg_6,data_in_shift_reg_5,data_in_shift_reg_4,data_in_shift_reg_3,data_in_shift_reg_2,data_in_shift_reg_1}),
	.comb(comb1),
	.GND_port(GND_port));

endmodule

module niosII_scfifo_5 (
	clock,
	q,
	full_dff,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	empty_dff,
	all_bits_transmitted,
	wrreq,
	data,
	comb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
output 	full_dff;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
output 	empty_dff;
input 	all_bits_transmitted;
input 	wrreq;
input 	[7:0] data;
input 	comb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_a341_2 auto_generated(
	.clock(clock),
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.full_dff(full_dff),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.all_bits_transmitted(all_bits_transmitted),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.comb(comb),
	.GND_port(GND_port));

endmodule

module niosII_scfifo_a341_2 (
	clock,
	q,
	full_dff,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	empty_dff,
	all_bits_transmitted,
	wrreq,
	data,
	comb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
output 	full_dff;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
output 	empty_dff;
input 	all_bits_transmitted;
input 	wrreq;
input 	[7:0] data;
input 	comb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_a_dpfifo_tq31_2 dpfifo(
	.clock(clock),
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.full_dff1(full_dff),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.r_sync_rst(r_sync_rst),
	.empty_dff1(empty_dff),
	.all_bits_transmitted(all_bits_transmitted),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.comb(comb),
	.GND_port(GND_port));

endmodule

module niosII_a_dpfifo_tq31_2 (
	clock,
	q,
	full_dff1,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	empty_dff1,
	all_bits_transmitted,
	wreq,
	data,
	comb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
output 	full_dff1;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
output 	empty_dff1;
input 	all_bits_transmitted;
input 	wreq;
input 	[7:0] data;
input 	comb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \wr_ptr|counter_reg_bit[6]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[5]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[5]~q ;
wire \ram_read_address[5]~5_combout ;
wire \low_addressa[6]~q ;
wire \ram_read_address[6]~6_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \low_addressa[5]~5_combout ;
wire \low_addressa[6]~6_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_will_be_1~4_combout ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \usedw_will_be_2~0_combout ;
wire \usedw_will_be_2~1_combout ;
wire \usedw_is_2_dff~q ;
wire \usedw_will_be_0~0_combout ;
wire \usedw_will_be_0~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~2_combout ;


niosII_cntr_0ab_2 wr_ptr(
	.clock(clock),
	.full_dff(full_dff1),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\wr_ptr|counter_reg_bit[6]~q ),
	.r_sync_rst(r_sync_rst),
	.all_bits_transmitted(all_bits_transmitted),
	.GND_port(GND_port));

niosII_cntr_ca7_2 usedw_counter(
	.clock(clock),
	.full_dff(full_dff1),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.r_sync_rst(r_sync_rst),
	.all_bits_transmitted(all_bits_transmitted),
	.updown(wreq),
	.comb(comb),
	.GND_port(GND_port));

niosII_cntr_v9b_2 rd_ptr_msb(
	.clock(clock),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.r_sync_rst(r_sync_rst),
	.comb(comb),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port));

niosII_altsyncram_dqb1_2 FIFOram(
	.clock0(clock),
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[6]~q ,\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_b({\ram_read_address[6]~6_combout ,\ram_read_address[5]~5_combout ,\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(comb),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

dffeas \low_addressa[5] (
	.clk(clock),
	.d(\low_addressa[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[5]~q ),
	.prn(vcc));
defparam \low_addressa[5] .is_wysiwyg = "true";
defparam \low_addressa[5] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[5]~5_combout ),
	.cout());
defparam \ram_read_address[5]~5 .lut_mask = 16'hAACC;
defparam \ram_read_address[5]~5 .sum_lutc_input = "datac";

dffeas \low_addressa[6] (
	.clk(clock),
	.d(\low_addressa[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[6]~q ),
	.prn(vcc));
defparam \low_addressa[6] .is_wysiwyg = "true";
defparam \low_addressa[6] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(gnd),
	.datad(comb),
	.cin(gnd),
	.combout(\ram_read_address[6]~6_combout ),
	.cout());
defparam \ram_read_address[6]~6 .lut_mask = 16'hAACC;
defparam \ram_read_address[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(comb),
	.datac(\rd_ptr_lsb~q ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'h8BFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(r_sync_rst),
	.datab(\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'h7777;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(r_sync_rst),
	.datab(comb),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEEEE;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hACFF;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hACFF;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hACFF;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hACFF;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[5]~5_combout ),
	.cout());
defparam \low_addressa[5]~5 .lut_mask = 16'hACFF;
defparam \low_addressa[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(comb),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[6]~6_combout ),
	.cout());
defparam \low_addressa[6]~6 .lut_mask = 16'hACFF;
defparam \low_addressa[6]~6 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \_~0 (
	.dataa(counter_reg_bit_6),
	.datab(counter_reg_bit_5),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_3),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFFE;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(all_bits_transmitted),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_2),
	.datad(\_~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(counter_reg_bit_1),
	.datab(full_dff1),
	.datac(comb),
	.datad(\_~1_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFFEF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~4 (
	.dataa(all_bits_transmitted),
	.datab(full_dff1),
	.datac(\usedw_is_1_dff~q ),
	.datad(comb),
	.cin(gnd),
	.combout(\usedw_will_be_1~4_combout ),
	.cout());
defparam \usedw_will_be_1~4 .lut_mask = 16'hF9F6;
defparam \usedw_will_be_1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_6),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hEFFF;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~4 (
	.dataa(\_~3_combout ),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_2),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hBFFF;
defparam \_~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~0 (
	.dataa(\_~4_combout ),
	.datab(\usedw_is_1_dff~q ),
	.datac(wreq),
	.datad(comb),
	.cin(gnd),
	.combout(\usedw_will_be_2~0_combout ),
	.cout());
defparam \usedw_will_be_2~0 .lut_mask = 16'hEFFE;
defparam \usedw_will_be_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~1 (
	.dataa(\usedw_will_be_2~0_combout ),
	.datab(\usedw_is_2_dff~q ),
	.datac(wreq),
	.datad(comb),
	.cin(gnd),
	.combout(\usedw_will_be_2~1_combout ),
	.cout());
defparam \usedw_will_be_2~1 .lut_mask = 16'hEFFE;
defparam \usedw_will_be_2~1 .sum_lutc_input = "datac";

dffeas usedw_is_2_dff(
	.clk(clock),
	.d(\usedw_will_be_2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_2_dff~q ),
	.prn(vcc));
defparam usedw_is_2_dff.is_wysiwyg = "true";
defparam usedw_is_2_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_0~0 (
	.dataa(wreq),
	.datab(comb),
	.datac(\usedw_is_1_dff~q ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\usedw_will_be_0~0_combout ),
	.cout());
defparam \usedw_will_be_0~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~1 (
	.dataa(\usedw_will_be_0~0_combout ),
	.datab(\usedw_is_0_dff~q ),
	.datac(wreq),
	.datad(comb),
	.cin(gnd),
	.combout(\usedw_will_be_0~1_combout ),
	.cout());
defparam \usedw_will_be_0~1 .lut_mask = 16'hEFFE;
defparam \usedw_will_be_0~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\usedw_will_be_0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(comb),
	.datac(\usedw_is_0_dff~q ),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFEF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(\usedw_will_be_1~4_combout ),
	.datab(\usedw_will_be_1~2_combout ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hEEFF;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(all_bits_transmitted),
	.datab(full_dff1),
	.datac(\usedw_will_be_1~3_combout ),
	.datad(\usedw_will_be_0~1_combout ),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hFFDF;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module niosII_altsyncram_dqb1_2 (
	clock0,
	q_b,
	address_a,
	wren_a,
	data_a,
	address_b)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[7:0] q_b;
input 	[6:0] address_a;
input 	wren_a;
input 	[7:0] data_a;
input 	[6:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_in_deserializer:RS232_In_Deserializer|altera_up_sync_fifo:RS232_In_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module niosII_cntr_0ab_2 (
	clock,
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	r_sync_rst,
	all_bits_transmitted,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	r_sync_rst;
input 	all_bits_transmitted;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(r_sync_rst),
	.datab(all_bits_transmitted),
	.datac(gnd),
	.datad(full_dff),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hEEFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module niosII_cntr_ca7_2 (
	clock,
	full_dff,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	r_sync_rst,
	all_bits_transmitted,
	updown,
	comb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	full_dff;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	r_sync_rst;
input 	all_bits_transmitted;
input 	updown;
input 	comb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;
wire \_~2_combout ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A6F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(all_bits_transmitted),
	.datab(full_dff),
	.datac(r_sync_rst),
	.datad(comb),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hF9F6;
defparam \_~2 .sum_lutc_input = "datac";

endmodule

module niosII_cntr_v9b_2 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	r_sync_rst,
	comb,
	rd_ptr_lsb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	r_sync_rst;
input 	comb;
input 	rd_ptr_lsb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(r_sync_rst),
	.datab(comb),
	.datac(gnd),
	.datad(rd_ptr_lsb),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hEEFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_altera_up_rs232_out_serializer_1 (
	wire_pll7_clk_0,
	write_fifo_write_en,
	fifo_write_space_7,
	fifo_write_space_6,
	fifo_write_space_5,
	fifo_write_space_4,
	fifo_write_space_3,
	fifo_write_space_2,
	fifo_write_space_1,
	fifo_write_space_0,
	serial_data_out1,
	r_sync_rst,
	data_to_uart_0,
	data_to_uart_1,
	data_to_uart_2,
	data_to_uart_3,
	data_to_uart_4,
	data_to_uart_5,
	data_to_uart_6,
	data_to_uart_7,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	write_fifo_write_en;
output 	fifo_write_space_7;
output 	fifo_write_space_6;
output 	fifo_write_space_5;
output 	fifo_write_space_4;
output 	fifo_write_space_3;
output 	fifo_write_space_2;
output 	fifo_write_space_1;
output 	fifo_write_space_0;
output 	serial_data_out1;
input 	r_sync_rst;
input 	data_to_uart_0;
input 	data_to_uart_1;
input 	data_to_uart_2;
input 	data_to_uart_3;
input 	data_to_uart_4;
input 	data_to_uart_5;
input 	data_to_uart_6;
input 	data_to_uart_7;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \RS232_Out_Counters|baud_clock_rising_edge~q ;
wire \RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \RS232_Out_Counters|all_bits_transmitted~q ;
wire \comb~0_combout ;
wire \data_out_shift_reg[6]~4_combout ;
wire \fifo_write_space[0]~9 ;
wire \fifo_write_space[1]~11 ;
wire \fifo_write_space[2]~13 ;
wire \fifo_write_space[3]~15 ;
wire \fifo_write_space[4]~17 ;
wire \fifo_write_space[5]~19 ;
wire \fifo_write_space[6]~21 ;
wire \fifo_write_space[7]~22_combout ;
wire \fifo_write_space[6]~20_combout ;
wire \fifo_write_space[5]~18_combout ;
wire \fifo_write_space[4]~16_combout ;
wire \fifo_write_space[3]~14_combout ;
wire \fifo_write_space[2]~12_combout ;
wire \fifo_write_space[1]~10_combout ;
wire \fifo_write_space[0]~8_combout ;
wire \transmitting_data~0_combout ;
wire \transmitting_data~q ;
wire \read_fifo_en~0_combout ;
wire \data_out_shift_reg~10_combout ;
wire \data_out_shift_reg[8]~q ;
wire \data_out_shift_reg~9_combout ;
wire \data_out_shift_reg[6]~2_combout ;
wire \data_out_shift_reg[7]~q ;
wire \data_out_shift_reg~8_combout ;
wire \data_out_shift_reg[6]~q ;
wire \data_out_shift_reg~7_combout ;
wire \data_out_shift_reg[5]~q ;
wire \data_out_shift_reg~6_combout ;
wire \data_out_shift_reg[4]~q ;
wire \data_out_shift_reg~5_combout ;
wire \data_out_shift_reg[3]~q ;
wire \data_out_shift_reg~3_combout ;
wire \data_out_shift_reg[2]~q ;
wire \data_out_shift_reg~1_combout ;
wire \data_out_shift_reg[1]~q ;
wire \data_out_shift_reg~0_combout ;
wire \data_out_shift_reg[0]~q ;
wire \serial_data_out~0_combout ;


niosII_altera_up_sync_fifo_3 RS232_Out_FIFO(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.q_b_0(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.q_b_1(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.counter_reg_bit_1(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_3(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_5(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_2(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_6(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.q_b_2(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.r_sync_rst(r_sync_rst),
	.empty_dff(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.read_fifo_en(\read_fifo_en~0_combout ),
	.comb(\comb~0_combout ),
	.data_to_uart_0(data_to_uart_0),
	.data_to_uart_1(data_to_uart_1),
	.data_out_shift_reg_6(\data_out_shift_reg[6]~4_combout ),
	.data_to_uart_2(data_to_uart_2),
	.data_to_uart_3(data_to_uart_3),
	.data_to_uart_4(data_to_uart_4),
	.data_to_uart_5(data_to_uart_5),
	.data_to_uart_6(data_to_uart_6),
	.data_to_uart_7(data_to_uart_7),
	.GND_port(GND_port));

niosII_altera_up_rs232_counters_3 RS232_Out_Counters(
	.clk(wire_pll7_clk_0),
	.transmitting_data(\transmitting_data~q ),
	.r_sync_rst(r_sync_rst),
	.baud_clock_rising_edge1(\RS232_Out_Counters|baud_clock_rising_edge~q ),
	.all_bits_transmitted1(\RS232_Out_Counters|all_bits_transmitted~q ));

cycloneive_lcell_comb \comb~0 (
	.dataa(write_fifo_write_en),
	.datab(gnd),
	.datac(gnd),
	.datad(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hAAFF;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg[6]~4 (
	.dataa(r_sync_rst),
	.datab(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datac(\RS232_Out_Counters|all_bits_transmitted~q ),
	.datad(\transmitting_data~q ),
	.cin(gnd),
	.combout(\data_out_shift_reg[6]~4_combout ),
	.cout());
defparam \data_out_shift_reg[6]~4 .lut_mask = 16'hEFFF;
defparam \data_out_shift_reg[6]~4 .sum_lutc_input = "datac";

dffeas \fifo_write_space[7] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_7),
	.prn(vcc));
defparam \fifo_write_space[7] .is_wysiwyg = "true";
defparam \fifo_write_space[7] .power_up = "low";

dffeas \fifo_write_space[6] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_6),
	.prn(vcc));
defparam \fifo_write_space[6] .is_wysiwyg = "true";
defparam \fifo_write_space[6] .power_up = "low";

dffeas \fifo_write_space[5] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_5),
	.prn(vcc));
defparam \fifo_write_space[5] .is_wysiwyg = "true";
defparam \fifo_write_space[5] .power_up = "low";

dffeas \fifo_write_space[4] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_4),
	.prn(vcc));
defparam \fifo_write_space[4] .is_wysiwyg = "true";
defparam \fifo_write_space[4] .power_up = "low";

dffeas \fifo_write_space[3] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_3),
	.prn(vcc));
defparam \fifo_write_space[3] .is_wysiwyg = "true";
defparam \fifo_write_space[3] .power_up = "low";

dffeas \fifo_write_space[2] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_2),
	.prn(vcc));
defparam \fifo_write_space[2] .is_wysiwyg = "true";
defparam \fifo_write_space[2] .power_up = "low";

dffeas \fifo_write_space[1] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_1),
	.prn(vcc));
defparam \fifo_write_space[1] .is_wysiwyg = "true";
defparam \fifo_write_space[1] .power_up = "low";

dffeas \fifo_write_space[0] (
	.clk(wire_pll7_clk_0),
	.d(\fifo_write_space[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_write_space_0),
	.prn(vcc));
defparam \fifo_write_space[0] .is_wysiwyg = "true";
defparam \fifo_write_space[0] .power_up = "low";

dffeas serial_data_out(
	.clk(wire_pll7_clk_0),
	.d(\serial_data_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(serial_data_out1),
	.prn(vcc));
defparam serial_data_out.is_wysiwyg = "true";
defparam serial_data_out.power_up = "low";

cycloneive_lcell_comb \fifo_write_space[0]~8 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\fifo_write_space[0]~8_combout ),
	.cout(\fifo_write_space[0]~9 ));
defparam \fifo_write_space[0]~8 .lut_mask = 16'hAA55;
defparam \fifo_write_space[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_write_space[1]~10 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[0]~9 ),
	.combout(\fifo_write_space[1]~10_combout ),
	.cout(\fifo_write_space[1]~11 ));
defparam \fifo_write_space[1]~10 .lut_mask = 16'h5AAF;
defparam \fifo_write_space[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[2]~12 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[1]~11 ),
	.combout(\fifo_write_space[2]~12_combout ),
	.cout(\fifo_write_space[2]~13 ));
defparam \fifo_write_space[2]~12 .lut_mask = 16'h5A5F;
defparam \fifo_write_space[2]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[3]~14 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[2]~13 ),
	.combout(\fifo_write_space[3]~14_combout ),
	.cout(\fifo_write_space[3]~15 ));
defparam \fifo_write_space[3]~14 .lut_mask = 16'h5AAF;
defparam \fifo_write_space[3]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[4]~16 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[3]~15 ),
	.combout(\fifo_write_space[4]~16_combout ),
	.cout(\fifo_write_space[4]~17 ));
defparam \fifo_write_space[4]~16 .lut_mask = 16'h5A5F;
defparam \fifo_write_space[4]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[5]~18 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[4]~17 ),
	.combout(\fifo_write_space[5]~18_combout ),
	.cout(\fifo_write_space[5]~19 ));
defparam \fifo_write_space[5]~18 .lut_mask = 16'h5AAF;
defparam \fifo_write_space[5]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[6]~20 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fifo_write_space[5]~19 ),
	.combout(\fifo_write_space[6]~20_combout ),
	.cout(\fifo_write_space[6]~21 ));
defparam \fifo_write_space[6]~20 .lut_mask = 16'h5A5F;
defparam \fifo_write_space[6]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fifo_write_space[7]~22 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fifo_write_space[6]~21 ),
	.combout(\fifo_write_space[7]~22_combout ),
	.cout());
defparam \fifo_write_space[7]~22 .lut_mask = 16'h5A5A;
defparam \fifo_write_space[7]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \transmitting_data~0 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datab(\transmitting_data~q ),
	.datac(gnd),
	.datad(\RS232_Out_Counters|all_bits_transmitted~q ),
	.cin(gnd),
	.combout(\transmitting_data~0_combout ),
	.cout());
defparam \transmitting_data~0 .lut_mask = 16'hEEFF;
defparam \transmitting_data~0 .sum_lutc_input = "datac";

dffeas transmitting_data(
	.clk(wire_pll7_clk_0),
	.d(\transmitting_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\transmitting_data~q ),
	.prn(vcc));
defparam transmitting_data.is_wysiwyg = "true";
defparam transmitting_data.power_up = "low";

cycloneive_lcell_comb \read_fifo_en~0 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datab(gnd),
	.datac(\RS232_Out_Counters|all_bits_transmitted~q ),
	.datad(\transmitting_data~q ),
	.cin(gnd),
	.combout(\read_fifo_en~0_combout ),
	.cout());
defparam \read_fifo_en~0 .lut_mask = 16'hAFFF;
defparam \read_fifo_en~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg~10 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(\RS232_Out_Counters|baud_clock_rising_edge~q ),
	.datac(\data_out_shift_reg[8]~q ),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~10_combout ),
	.cout());
defparam \data_out_shift_reg~10 .lut_mask = 16'hFAFC;
defparam \data_out_shift_reg~10 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[8] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(vcc),
	.q(\data_out_shift_reg[8]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[8] .is_wysiwyg = "true";
defparam \data_out_shift_reg[8] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~9 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(\data_out_shift_reg[8]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~9_combout ),
	.cout());
defparam \data_out_shift_reg~9 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg[6]~2 (
	.dataa(r_sync_rst),
	.datab(\RS232_Out_Counters|baud_clock_rising_edge~q ),
	.datac(\read_fifo_en~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_out_shift_reg[6]~2_combout ),
	.cout());
defparam \data_out_shift_reg[6]~2 .lut_mask = 16'hFEFE;
defparam \data_out_shift_reg[6]~2 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[7] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[6]~2_combout ),
	.q(\data_out_shift_reg[7]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[7] .is_wysiwyg = "true";
defparam \data_out_shift_reg[7] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~8 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(\data_out_shift_reg[7]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~8_combout ),
	.cout());
defparam \data_out_shift_reg~8 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~8 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[6] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[6]~2_combout ),
	.q(\data_out_shift_reg[6]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[6] .is_wysiwyg = "true";
defparam \data_out_shift_reg[6] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~7 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datab(\data_out_shift_reg[6]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~7_combout ),
	.cout());
defparam \data_out_shift_reg~7 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~7 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[5] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[6]~2_combout ),
	.q(\data_out_shift_reg[5]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[5] .is_wysiwyg = "true";
defparam \data_out_shift_reg[5] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~6 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datab(\data_out_shift_reg[5]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~6_combout ),
	.cout());
defparam \data_out_shift_reg~6 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~6 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[4] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[6]~2_combout ),
	.q(\data_out_shift_reg[4]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[4] .is_wysiwyg = "true";
defparam \data_out_shift_reg[4] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~5 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(\data_out_shift_reg[4]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~5_combout ),
	.cout());
defparam \data_out_shift_reg~5 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~5 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[3] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[6]~2_combout ),
	.q(\data_out_shift_reg[3]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[3] .is_wysiwyg = "true";
defparam \data_out_shift_reg[3] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~3 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(\data_out_shift_reg[3]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~3_combout ),
	.cout());
defparam \data_out_shift_reg~3 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~3 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[2] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[6]~2_combout ),
	.q(\data_out_shift_reg[2]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[2] .is_wysiwyg = "true";
defparam \data_out_shift_reg[2] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~1 (
	.dataa(\RS232_Out_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\data_out_shift_reg[2]~q ),
	.datac(gnd),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~1_combout ),
	.cout());
defparam \data_out_shift_reg~1 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg~1 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[1] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\data_out_shift_reg[6]~2_combout ),
	.q(\data_out_shift_reg[1]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[1] .is_wysiwyg = "true";
defparam \data_out_shift_reg[1] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg~0 (
	.dataa(\data_out_shift_reg[1]~q ),
	.datab(\data_out_shift_reg[0]~q ),
	.datac(\RS232_Out_Counters|baud_clock_rising_edge~q ),
	.datad(\read_fifo_en~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~0_combout ),
	.cout());
defparam \data_out_shift_reg~0 .lut_mask = 16'hACFF;
defparam \data_out_shift_reg~0 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[0] (
	.clk(wire_pll7_clk_0),
	.d(\data_out_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(vcc),
	.q(\data_out_shift_reg[0]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[0] .is_wysiwyg = "true";
defparam \data_out_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \serial_data_out~0 (
	.dataa(r_sync_rst),
	.datab(\data_out_shift_reg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\serial_data_out~0_combout ),
	.cout());
defparam \serial_data_out~0 .lut_mask = 16'hEEEE;
defparam \serial_data_out~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_rs232_counters_3 (
	clk,
	transmitting_data,
	r_sync_rst,
	baud_clock_rising_edge1,
	all_bits_transmitted1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	transmitting_data;
input 	r_sync_rst;
output 	baud_clock_rising_edge1;
output 	all_bits_transmitted1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \baud_counter[0]~10_combout ;
wire \baud_counter[9]~12_combout ;
wire \baud_counter[0]~q ;
wire \baud_counter[0]~11 ;
wire \baud_counter[1]~13_combout ;
wire \baud_counter[1]~q ;
wire \baud_counter[1]~14 ;
wire \baud_counter[2]~15_combout ;
wire \baud_counter[2]~q ;
wire \baud_counter[2]~16 ;
wire \baud_counter[3]~17_combout ;
wire \baud_counter[3]~q ;
wire \Equal0~0_combout ;
wire \baud_counter[3]~18 ;
wire \baud_counter[4]~19_combout ;
wire \baud_counter[4]~q ;
wire \baud_counter[4]~20 ;
wire \baud_counter[5]~21_combout ;
wire \baud_counter[5]~q ;
wire \baud_counter[5]~22 ;
wire \baud_counter[6]~23_combout ;
wire \baud_counter[6]~q ;
wire \baud_counter[6]~24 ;
wire \baud_counter[7]~25_combout ;
wire \baud_counter[7]~q ;
wire \Equal0~1_combout ;
wire \baud_counter[7]~26 ;
wire \baud_counter[8]~27_combout ;
wire \baud_counter[8]~q ;
wire \baud_counter[8]~28 ;
wire \baud_counter[9]~29_combout ;
wire \baud_counter[9]~q ;
wire \Equal0~2_combout ;
wire \baud_clock_rising_edge~0_combout ;
wire \bit_counter[2]~0_combout ;
wire \bit_counter[0]~2_combout ;
wire \bit_counter[0]~q ;
wire \bit_counter[1]~3_combout ;
wire \bit_counter[1]~q ;
wire \Add1~0_combout ;
wire \bit_counter[2]~1_combout ;
wire \bit_counter[2]~q ;
wire \Add1~1_combout ;
wire \bit_counter[3]~4_combout ;
wire \bit_counter[3]~q ;
wire \Equal2~0_combout ;
wire \all_bits_transmitted~0_combout ;


dffeas baud_clock_rising_edge(
	.clk(clk),
	.d(\baud_clock_rising_edge~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(baud_clock_rising_edge1),
	.prn(vcc));
defparam baud_clock_rising_edge.is_wysiwyg = "true";
defparam baud_clock_rising_edge.power_up = "low";

dffeas all_bits_transmitted(
	.clk(clk),
	.d(\all_bits_transmitted~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(all_bits_transmitted1),
	.prn(vcc));
defparam all_bits_transmitted.is_wysiwyg = "true";
defparam all_bits_transmitted.power_up = "low";

cycloneive_lcell_comb \baud_counter[0]~10 (
	.dataa(\baud_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\baud_counter[0]~10_combout ),
	.cout(\baud_counter[0]~11 ));
defparam \baud_counter[0]~10 .lut_mask = 16'h55AA;
defparam \baud_counter[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[9]~12 (
	.dataa(transmitting_data),
	.datab(\Equal0~2_combout ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\baud_counter[9]~12_combout ),
	.cout());
defparam \baud_counter[9]~12 .lut_mask = 16'hFF77;
defparam \baud_counter[9]~12 .sum_lutc_input = "datac";

dffeas \baud_counter[0] (
	.clk(clk),
	.d(\baud_counter[0]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[0]~q ),
	.prn(vcc));
defparam \baud_counter[0] .is_wysiwyg = "true";
defparam \baud_counter[0] .power_up = "low";

cycloneive_lcell_comb \baud_counter[1]~13 (
	.dataa(\baud_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[0]~11 ),
	.combout(\baud_counter[1]~13_combout ),
	.cout(\baud_counter[1]~14 ));
defparam \baud_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \baud_counter[1]~13 .sum_lutc_input = "cin";

dffeas \baud_counter[1] (
	.clk(clk),
	.d(\baud_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[1]~q ),
	.prn(vcc));
defparam \baud_counter[1] .is_wysiwyg = "true";
defparam \baud_counter[1] .power_up = "low";

cycloneive_lcell_comb \baud_counter[2]~15 (
	.dataa(\baud_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[1]~14 ),
	.combout(\baud_counter[2]~15_combout ),
	.cout(\baud_counter[2]~16 ));
defparam \baud_counter[2]~15 .lut_mask = 16'h5AAF;
defparam \baud_counter[2]~15 .sum_lutc_input = "cin";

dffeas \baud_counter[2] (
	.clk(clk),
	.d(\baud_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[2]~q ),
	.prn(vcc));
defparam \baud_counter[2] .is_wysiwyg = "true";
defparam \baud_counter[2] .power_up = "low";

cycloneive_lcell_comb \baud_counter[3]~17 (
	.dataa(\baud_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[2]~16 ),
	.combout(\baud_counter[3]~17_combout ),
	.cout(\baud_counter[3]~18 ));
defparam \baud_counter[3]~17 .lut_mask = 16'h5A5F;
defparam \baud_counter[3]~17 .sum_lutc_input = "cin";

dffeas \baud_counter[3] (
	.clk(clk),
	.d(\baud_counter[3]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[3]~q ),
	.prn(vcc));
defparam \baud_counter[3] .is_wysiwyg = "true";
defparam \baud_counter[3] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\baud_counter[0]~q ),
	.datab(\baud_counter[1]~q ),
	.datac(\baud_counter[3]~q ),
	.datad(\baud_counter[2]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFEFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[4]~19 (
	.dataa(\baud_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[3]~18 ),
	.combout(\baud_counter[4]~19_combout ),
	.cout(\baud_counter[4]~20 ));
defparam \baud_counter[4]~19 .lut_mask = 16'h5AAF;
defparam \baud_counter[4]~19 .sum_lutc_input = "cin";

dffeas \baud_counter[4] (
	.clk(clk),
	.d(\baud_counter[4]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[4]~q ),
	.prn(vcc));
defparam \baud_counter[4] .is_wysiwyg = "true";
defparam \baud_counter[4] .power_up = "low";

cycloneive_lcell_comb \baud_counter[5]~21 (
	.dataa(\baud_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[4]~20 ),
	.combout(\baud_counter[5]~21_combout ),
	.cout(\baud_counter[5]~22 ));
defparam \baud_counter[5]~21 .lut_mask = 16'h5A5F;
defparam \baud_counter[5]~21 .sum_lutc_input = "cin";

dffeas \baud_counter[5] (
	.clk(clk),
	.d(\baud_counter[5]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[5]~q ),
	.prn(vcc));
defparam \baud_counter[5] .is_wysiwyg = "true";
defparam \baud_counter[5] .power_up = "low";

cycloneive_lcell_comb \baud_counter[6]~23 (
	.dataa(\baud_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[5]~22 ),
	.combout(\baud_counter[6]~23_combout ),
	.cout(\baud_counter[6]~24 ));
defparam \baud_counter[6]~23 .lut_mask = 16'h5AAF;
defparam \baud_counter[6]~23 .sum_lutc_input = "cin";

dffeas \baud_counter[6] (
	.clk(clk),
	.d(\baud_counter[6]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[6]~q ),
	.prn(vcc));
defparam \baud_counter[6] .is_wysiwyg = "true";
defparam \baud_counter[6] .power_up = "low";

cycloneive_lcell_comb \baud_counter[7]~25 (
	.dataa(\baud_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[6]~24 ),
	.combout(\baud_counter[7]~25_combout ),
	.cout(\baud_counter[7]~26 ));
defparam \baud_counter[7]~25 .lut_mask = 16'h5A5F;
defparam \baud_counter[7]~25 .sum_lutc_input = "cin";

dffeas \baud_counter[7] (
	.clk(clk),
	.d(\baud_counter[7]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[7]~q ),
	.prn(vcc));
defparam \baud_counter[7] .is_wysiwyg = "true";
defparam \baud_counter[7] .power_up = "low";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\baud_counter[4]~q ),
	.datab(\baud_counter[7]~q ),
	.datac(\baud_counter[5]~q ),
	.datad(\baud_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_counter[8]~27 (
	.dataa(\baud_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\baud_counter[7]~26 ),
	.combout(\baud_counter[8]~27_combout ),
	.cout(\baud_counter[8]~28 ));
defparam \baud_counter[8]~27 .lut_mask = 16'h5AAF;
defparam \baud_counter[8]~27 .sum_lutc_input = "cin";

dffeas \baud_counter[8] (
	.clk(clk),
	.d(\baud_counter[8]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[8]~q ),
	.prn(vcc));
defparam \baud_counter[8] .is_wysiwyg = "true";
defparam \baud_counter[8] .power_up = "low";

cycloneive_lcell_comb \baud_counter[9]~29 (
	.dataa(\baud_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\baud_counter[8]~28 ),
	.combout(\baud_counter[9]~29_combout ),
	.cout());
defparam \baud_counter[9]~29 .lut_mask = 16'h5A5A;
defparam \baud_counter[9]~29 .sum_lutc_input = "cin";

dffeas \baud_counter[9] (
	.clk(clk),
	.d(\baud_counter[9]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\baud_counter[9]~12_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\baud_counter[9]~q ),
	.prn(vcc));
defparam \baud_counter[9] .is_wysiwyg = "true";
defparam \baud_counter[9] .power_up = "low";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\baud_counter[8]~q ),
	.datad(\baud_counter[9]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEFFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \baud_clock_rising_edge~0 (
	.dataa(r_sync_rst),
	.datab(\Equal0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\baud_clock_rising_edge~0_combout ),
	.cout());
defparam \baud_clock_rising_edge~0 .lut_mask = 16'h7777;
defparam \baud_clock_rising_edge~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[2]~0 (
	.dataa(transmitting_data),
	.datab(\Equal2~0_combout ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\bit_counter[2]~0_combout ),
	.cout());
defparam \bit_counter[2]~0 .lut_mask = 16'hEEFF;
defparam \bit_counter[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[0]~2 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\Equal0~2_combout ),
	.datac(\bit_counter[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\bit_counter[0]~2_combout ),
	.cout());
defparam \bit_counter[0]~2 .lut_mask = 16'hBEBE;
defparam \bit_counter[0]~2 .sum_lutc_input = "datac";

dffeas \bit_counter[0] (
	.clk(clk),
	.d(\bit_counter[0]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[0]~q ),
	.prn(vcc));
defparam \bit_counter[0] .is_wysiwyg = "true";
defparam \bit_counter[0] .power_up = "low";

cycloneive_lcell_comb \bit_counter[1]~3 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[1]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\bit_counter[1]~3_combout ),
	.cout());
defparam \bit_counter[1]~3 .lut_mask = 16'hEBBE;
defparam \bit_counter[1]~3 .sum_lutc_input = "datac";

dffeas \bit_counter[1] (
	.clk(clk),
	.d(\bit_counter[1]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[1]~q ),
	.prn(vcc));
defparam \bit_counter[1] .is_wysiwyg = "true";
defparam \bit_counter[1] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(\bit_counter[2]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'hC33C;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[2]~1 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[2]~q ),
	.datac(\Add1~0_combout ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\bit_counter[2]~1_combout ),
	.cout());
defparam \bit_counter[2]~1 .lut_mask = 16'hFAFC;
defparam \bit_counter[2]~1 .sum_lutc_input = "datac";

dffeas \bit_counter[2] (
	.clk(clk),
	.d(\bit_counter[2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[2]~q ),
	.prn(vcc));
defparam \bit_counter[2] .is_wysiwyg = "true";
defparam \bit_counter[2] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(\bit_counter[3]~q ),
	.datab(\bit_counter[2]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[0]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[3]~4 (
	.dataa(\bit_counter[2]~0_combout ),
	.datab(\bit_counter[3]~q ),
	.datac(\Add1~1_combout ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\bit_counter[3]~4_combout ),
	.cout());
defparam \bit_counter[3]~4 .lut_mask = 16'hFAFC;
defparam \bit_counter[3]~4 .sum_lutc_input = "datac";

dffeas \bit_counter[3] (
	.clk(clk),
	.d(\bit_counter[3]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_counter[3]~q ),
	.prn(vcc));
defparam \bit_counter[3] .is_wysiwyg = "true";
defparam \bit_counter[3] .power_up = "low";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(\bit_counter[2]~q ),
	.datab(\bit_counter[0]~q ),
	.datac(\bit_counter[1]~q ),
	.datad(\bit_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hEFFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \all_bits_transmitted~0 (
	.dataa(r_sync_rst),
	.datab(\Equal2~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\all_bits_transmitted~0_combout ),
	.cout());
defparam \all_bits_transmitted~0 .lut_mask = 16'h7777;
defparam \all_bits_transmitted~0 .sum_lutc_input = "datac";

endmodule

module niosII_altera_up_sync_fifo_3 (
	wire_pll7_clk_0,
	q_b_0,
	write_fifo_write_en,
	full_dff,
	q_b_1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_2,
	counter_reg_bit_6,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	r_sync_rst,
	empty_dff,
	read_fifo_en,
	comb,
	data_to_uart_0,
	data_to_uart_1,
	data_out_shift_reg_6,
	data_to_uart_2,
	data_to_uart_3,
	data_to_uart_4,
	data_to_uart_5,
	data_to_uart_6,
	data_to_uart_7,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	q_b_0;
input 	write_fifo_write_en;
output 	full_dff;
output 	q_b_1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_2;
output 	counter_reg_bit_6;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	r_sync_rst;
output 	empty_dff;
input 	read_fifo_en;
input 	comb;
input 	data_to_uart_0;
input 	data_to_uart_1;
input 	data_out_shift_reg_6;
input 	data_to_uart_2;
input 	data_to_uart_3;
input 	data_to_uart_4;
input 	data_to_uart_5;
input 	data_to_uart_6;
input 	data_to_uart_7;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_6 Sync_FIFO(
	.clock(wire_pll7_clk_0),
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(full_dff),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_6(counter_reg_bit_6),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.read_fifo_en(read_fifo_en),
	.wrreq(comb),
	.data({data_to_uart_7,data_to_uart_6,data_to_uart_5,data_to_uart_4,data_to_uart_3,data_to_uart_2,data_to_uart_1,data_to_uart_0}),
	.data_out_shift_reg_6(data_out_shift_reg_6),
	.GND_port(GND_port));

endmodule

module niosII_scfifo_6 (
	clock,
	q,
	write_fifo_write_en,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_2,
	counter_reg_bit_6,
	r_sync_rst,
	empty_dff,
	read_fifo_en,
	wrreq,
	data,
	data_out_shift_reg_6,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
input 	write_fifo_write_en;
output 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_2;
output 	counter_reg_bit_6;
input 	r_sync_rst;
output 	empty_dff;
input 	read_fifo_en;
input 	wrreq;
input 	[7:0] data;
input 	data_out_shift_reg_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_scfifo_a341_3 auto_generated(
	.clock(clock),
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(full_dff),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_6(counter_reg_bit_6),
	.r_sync_rst(r_sync_rst),
	.empty_dff(empty_dff),
	.read_fifo_en(read_fifo_en),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.data_out_shift_reg_6(data_out_shift_reg_6),
	.GND_port(GND_port));

endmodule

module niosII_scfifo_a341_3 (
	clock,
	q,
	write_fifo_write_en,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_2,
	counter_reg_bit_6,
	r_sync_rst,
	empty_dff,
	read_fifo_en,
	wrreq,
	data,
	data_out_shift_reg_6,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
input 	write_fifo_write_en;
output 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_2;
output 	counter_reg_bit_6;
input 	r_sync_rst;
output 	empty_dff;
input 	read_fifo_en;
input 	wrreq;
input 	[7:0] data;
input 	data_out_shift_reg_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_a_dpfifo_tq31_3 dpfifo(
	.clock(clock),
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff1(full_dff),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_6(counter_reg_bit_6),
	.r_sync_rst(r_sync_rst),
	.empty_dff1(empty_dff),
	.read_fifo_en(read_fifo_en),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.data_out_shift_reg_6(data_out_shift_reg_6),
	.GND_port(GND_port));

endmodule

module niosII_a_dpfifo_tq31_3 (
	clock,
	q,
	write_fifo_write_en,
	full_dff1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_2,
	counter_reg_bit_6,
	r_sync_rst,
	empty_dff1,
	read_fifo_en,
	wreq,
	data,
	data_out_shift_reg_6,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[7:0] q;
input 	write_fifo_write_en;
output 	full_dff1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_2;
output 	counter_reg_bit_6;
input 	r_sync_rst;
output 	empty_dff1;
input 	read_fifo_en;
input 	wreq;
input 	[7:0] data;
input 	data_out_shift_reg_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \wr_ptr|counter_reg_bit[6]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[5]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[5]~q ;
wire \ram_read_address[5]~5_combout ;
wire \low_addressa[6]~q ;
wire \ram_read_address[6]~6_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \low_addressa[5]~5_combout ;
wire \low_addressa[6]~6_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_will_be_2~0_combout ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \usedw_will_be_2~1_combout ;
wire \usedw_is_2_dff~q ;
wire \usedw_will_be_1~4_combout ;
wire \usedw_will_be_0~0_combout ;
wire \usedw_will_be_0~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~0_combout ;


niosII_cntr_0ab_3 wr_ptr(
	.clock(clock),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(full_dff1),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\wr_ptr|counter_reg_bit[6]~q ),
	.r_sync_rst(r_sync_rst),
	.GND_port(GND_port));

niosII_cntr_ca7_3 usedw_counter(
	.clock(clock),
	.write_fifo_write_en(write_fifo_write_en),
	.full_dff(full_dff1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_6(counter_reg_bit_6),
	.r_sync_rst(r_sync_rst),
	.read_fifo_en(read_fifo_en),
	.updown(wreq),
	.GND_port(GND_port));

niosII_cntr_v9b_3 rd_ptr_msb(
	.clock(clock),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.r_sync_rst(r_sync_rst),
	.read_fifo_en(read_fifo_en),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port));

niosII_altsyncram_dqb1_3 FIFOram(
	.clock0(clock),
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[6]~q ,\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_b({\ram_read_address[6]~6_combout ,\ram_read_address[5]~5_combout ,\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_shift_reg_6),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(read_fifo_en),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

dffeas \low_addressa[5] (
	.clk(clock),
	.d(\low_addressa[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[5]~q ),
	.prn(vcc));
defparam \low_addressa[5] .is_wysiwyg = "true";
defparam \low_addressa[5] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[5]~5_combout ),
	.cout());
defparam \ram_read_address[5]~5 .lut_mask = 16'hAACC;
defparam \ram_read_address[5]~5 .sum_lutc_input = "datac";

dffeas \low_addressa[6] (
	.clk(clock),
	.d(\low_addressa[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[6]~q ),
	.prn(vcc));
defparam \low_addressa[6] .is_wysiwyg = "true";
defparam \low_addressa[6] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(gnd),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\ram_read_address[6]~6_combout ),
	.cout());
defparam \ram_read_address[6]~6 .lut_mask = 16'hAACC;
defparam \ram_read_address[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(read_fifo_en),
	.datac(\rd_ptr_lsb~q ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'h8BFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(r_sync_rst),
	.datab(\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'h7777;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hACFF;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hACFF;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hACFF;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hACFF;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[5]~5_combout ),
	.cout());
defparam \low_addressa[5]~5 .lut_mask = 16'hACFF;
defparam \low_addressa[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(read_fifo_en),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\low_addressa[6]~6_combout ),
	.cout());
defparam \low_addressa[6]~6 .lut_mask = 16'hACFF;
defparam \low_addressa[6]~6 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \_~0 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFFE;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(write_fifo_write_en),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_6),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(full_dff1),
	.datab(read_fifo_en),
	.datac(\_~0_combout ),
	.datad(\_~1_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFFFB;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_2~0 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\usedw_will_be_2~0_combout ),
	.cout());
defparam \usedw_will_be_2~0 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_6),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hEFFF;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~4 (
	.dataa(\_~3_combout ),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_3),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hBFFF;
defparam \_~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~1 (
	.dataa(\usedw_will_be_2~0_combout ),
	.datab(read_fifo_en),
	.datac(\_~4_combout ),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_2~1_combout ),
	.cout());
defparam \usedw_will_be_2~1 .lut_mask = 16'hFEFF;
defparam \usedw_will_be_2~1 .sum_lutc_input = "datac";

dffeas usedw_is_2_dff(
	.clk(clock),
	.d(\usedw_will_be_2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(r_sync_rst),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_2_dff~q ),
	.prn(vcc));
defparam usedw_is_2_dff.is_wysiwyg = "true";
defparam usedw_is_2_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~4 (
	.dataa(write_fifo_write_en),
	.datab(full_dff1),
	.datac(read_fifo_en),
	.datad(\usedw_is_2_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~4_combout ),
	.cout());
defparam \usedw_will_be_1~4 .lut_mask = 16'hFFFD;
defparam \usedw_will_be_1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\usedw_will_be_0~0_combout ),
	.cout());
defparam \usedw_will_be_0~0 .lut_mask = 16'hBFEF;
defparam \usedw_will_be_0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~1 (
	.dataa(\usedw_will_be_0~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\usedw_will_be_0~1_combout ),
	.cout());
defparam \usedw_will_be_0~1 .lut_mask = 16'hAAFF;
defparam \usedw_will_be_0~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\usedw_will_be_0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(wreq),
	.datac(read_fifo_en),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBEFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(\usedw_will_be_1~4_combout ),
	.datab(\usedw_will_be_1~2_combout ),
	.datac(gnd),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hEEFF;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(r_sync_rst),
	.datab(wreq),
	.datac(\usedw_will_be_1~3_combout ),
	.datad(\usedw_will_be_0~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hFF7F;
defparam \empty_dff~0 .sum_lutc_input = "datac";

endmodule

module niosII_altsyncram_dqb1_3 (
	clock0,
	q_b,
	address_a,
	wren_a,
	data_a,
	address_b)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[7:0] q_b;
input 	[6:0] address_a;
input 	wren_a;
input 	[7:0] data_a;
input 	[6:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosII_rs232_0:rs232_1|altera_up_rs232_out_serializer:RS232_Out_Serializer|altera_up_sync_fifo:RS232_Out_FIFO|scfifo:Sync_FIFO|scfifo_a341:auto_generated|a_dpfifo_tq31:dpfifo|altsyncram_dqb1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module niosII_cntr_0ab_3 (
	clock,
	write_fifo_write_en,
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	r_sync_rst,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	write_fifo_write_en;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	r_sync_rst;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(r_sync_rst),
	.datab(write_fifo_write_en),
	.datac(gnd),
	.datad(full_dff),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hEEFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module niosII_cntr_ca7_3 (
	clock,
	write_fifo_write_en,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_2,
	counter_reg_bit_6,
	r_sync_rst,
	read_fifo_en,
	updown,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	write_fifo_write_en;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_2;
output 	counter_reg_bit_6;
input 	r_sync_rst;
input 	read_fifo_en;
input 	updown;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(write_fifo_write_en),
	.datab(full_dff),
	.datac(r_sync_rst),
	.datad(read_fifo_en),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hF9F6;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A6F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module niosII_cntr_v9b_3 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	r_sync_rst,
	read_fifo_en,
	rd_ptr_lsb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	r_sync_rst;
input 	read_fifo_en;
input 	rd_ptr_lsb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(r_sync_rst),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(r_sync_rst),
	.datab(read_fifo_en),
	.datac(gnd),
	.datad(rd_ptr_lsb),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hEEFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module niosII_niosII_sdram (
	wire_pll7_clk_0,
	m_addr_0,
	m_addr_1,
	m_addr_2,
	m_addr_3,
	m_addr_4,
	m_addr_5,
	m_addr_6,
	m_addr_7,
	m_addr_8,
	byteen_reg_0,
	byteen_reg_1,
	oe1,
	m_addr_9,
	m_addr_10,
	m_addr_11,
	m_addr_12,
	m_bank_0,
	m_bank_1,
	m_cmd_1,
	m_cmd_3,
	m_dqm_0,
	m_dqm_1,
	m_cmd_2,
	m_cmd_0,
	r_sync_rst,
	entries_1,
	entries_0,
	d_byteenable_0,
	saved_grant_0,
	d_byteenable_1,
	use_reg,
	saved_grant_1,
	WideOr0,
	Equal0,
	Equal1,
	WideOr1,
	m0_write,
	mem_used_7,
	src_data_66,
	out_data_28,
	src_valid,
	src12_valid,
	m0_write1,
	out_data_42,
	out_data_29,
	out_data_31,
	out_data_30,
	out_data_33,
	out_data_32,
	out_data_35,
	out_data_34,
	out_data_37,
	out_data_36,
	out_data_39,
	out_data_38,
	out_data_41,
	out_data_40,
	out_data_19,
	out_data_20,
	out_data_21,
	out_data_22,
	out_data_23,
	out_data_24,
	out_data_25,
	out_data_26,
	out_data_27,
	m_data_0,
	m_data_1,
	m_data_2,
	m_data_3,
	m_data_4,
	m_data_5,
	m_data_6,
	m_data_7,
	m_data_8,
	m_data_9,
	m_data_10,
	m_data_11,
	m_data_12,
	m_data_13,
	m_data_14,
	m_data_15,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	za_valid1,
	za_data_0,
	za_data_1,
	za_data_2,
	za_data_3,
	za_data_4,
	za_data_11,
	za_data_13,
	za_data_12,
	za_data_5,
	za_data_14,
	za_data_15,
	za_data_10,
	za_data_9,
	za_data_8,
	za_data_7,
	za_data_6,
	sdram_dq_0,
	sdram_dq_1,
	sdram_dq_2,
	sdram_dq_3,
	sdram_dq_4,
	sdram_dq_5,
	sdram_dq_6,
	sdram_dq_7,
	sdram_dq_8,
	sdram_dq_9,
	sdram_dq_10,
	sdram_dq_11,
	sdram_dq_12,
	sdram_dq_13,
	sdram_dq_14,
	sdram_dq_15)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	m_addr_0;
output 	m_addr_1;
output 	m_addr_2;
output 	m_addr_3;
output 	m_addr_4;
output 	m_addr_5;
output 	m_addr_6;
output 	m_addr_7;
output 	m_addr_8;
input 	byteen_reg_0;
input 	byteen_reg_1;
output 	oe1;
output 	m_addr_9;
output 	m_addr_10;
output 	m_addr_11;
output 	m_addr_12;
output 	m_bank_0;
output 	m_bank_1;
output 	m_cmd_1;
output 	m_cmd_3;
output 	m_dqm_0;
output 	m_dqm_1;
output 	m_cmd_2;
output 	m_cmd_0;
input 	r_sync_rst;
output 	entries_1;
output 	entries_0;
input 	d_byteenable_0;
input 	saved_grant_0;
input 	d_byteenable_1;
input 	use_reg;
input 	saved_grant_1;
input 	WideOr0;
output 	Equal0;
input 	Equal1;
input 	WideOr1;
input 	m0_write;
input 	mem_used_7;
input 	src_data_66;
input 	out_data_28;
input 	src_valid;
input 	src12_valid;
input 	m0_write1;
input 	out_data_42;
input 	out_data_29;
input 	out_data_31;
input 	out_data_30;
input 	out_data_33;
input 	out_data_32;
input 	out_data_35;
input 	out_data_34;
input 	out_data_37;
input 	out_data_36;
input 	out_data_39;
input 	out_data_38;
input 	out_data_41;
input 	out_data_40;
input 	out_data_19;
input 	out_data_20;
input 	out_data_21;
input 	out_data_22;
input 	out_data_23;
input 	out_data_24;
input 	out_data_25;
input 	out_data_26;
input 	out_data_27;
output 	m_data_0;
output 	m_data_1;
output 	m_data_2;
output 	m_data_3;
output 	m_data_4;
output 	m_data_5;
output 	m_data_6;
output 	m_data_7;
output 	m_data_8;
output 	m_data_9;
output 	m_data_10;
output 	m_data_11;
output 	m_data_12;
output 	m_data_13;
output 	m_data_14;
output 	m_data_15;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
input 	out_data_5;
input 	out_data_6;
input 	out_data_7;
input 	out_data_8;
input 	out_data_9;
input 	out_data_10;
input 	out_data_11;
input 	out_data_12;
input 	out_data_13;
input 	out_data_14;
input 	out_data_15;
output 	za_valid1;
output 	za_data_0;
output 	za_data_1;
output 	za_data_2;
output 	za_data_3;
output 	za_data_4;
output 	za_data_11;
output 	za_data_13;
output 	za_data_12;
output 	za_data_5;
output 	za_data_14;
output 	za_data_15;
output 	za_data_10;
output 	za_data_9;
output 	za_data_8;
output 	za_data_7;
output 	za_data_6;
input 	sdram_dq_0;
input 	sdram_dq_1;
input 	sdram_dq_2;
input 	sdram_dq_3;
input 	sdram_dq_4;
input 	sdram_dq_5;
input 	sdram_dq_6;
input 	sdram_dq_7;
input 	sdram_dq_8;
input 	sdram_dq_9;
input 	sdram_dq_10;
input 	sdram_dq_11;
input 	sdram_dq_12;
input 	sdram_dq_13;
input 	sdram_dq_14;
input 	sdram_dq_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_niosII_sdram_input_efifo_module|Equal1~0_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[27]~0_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[42]~1_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[41]~2_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[28]~3_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[30]~4_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[29]~5_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[32]~6_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[31]~7_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[34]~8_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[33]~9_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[36]~10_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[35]~11_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[38]~12_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[37]~13_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[40]~14_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[39]~15_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[18]~16_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[19]~17_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[20]~18_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[21]~19_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[22]~20_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[23]~21_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[24]~22_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[25]~23_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[26]~24_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[16]~25_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[17]~26_combout ;
wire \comb~0_combout ;
wire \comb~1_combout ;
wire \comb~2_combout ;
wire \comb~3_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[0]~27_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[1]~28_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[2]~29_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[3]~30_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[4]~31_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[5]~32_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[6]~33_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[7]~34_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[8]~35_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[9]~36_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[10]~37_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[11]~38_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[12]~39_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[13]~40_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[14]~41_combout ;
wire \the_niosII_sdram_input_efifo_module|rd_data[15]~42_combout ;
wire \Add0~0_combout ;
wire \refresh_counter~8_combout ;
wire \refresh_counter[0]~q ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \refresh_counter[1]~q ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \refresh_counter~7_combout ;
wire \refresh_counter[2]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \refresh_counter[3]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \refresh_counter[4]~13_combout ;
wire \refresh_counter[4]~q ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \refresh_counter~6_combout ;
wire \refresh_counter[5]~q ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \refresh_counter~5_combout ;
wire \refresh_counter[6]~q ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \refresh_counter~4_combout ;
wire \refresh_counter[7]~q ;
wire \Add0~15 ;
wire \Add0~16_combout ;
wire \refresh_counter~3_combout ;
wire \refresh_counter[8]~q ;
wire \Add0~17 ;
wire \Add0~18_combout ;
wire \refresh_counter[9]~11_combout ;
wire \refresh_counter[9]~q ;
wire \Add0~19 ;
wire \Add0~20_combout ;
wire \refresh_counter[10]~10_combout ;
wire \refresh_counter[10]~q ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \refresh_counter~2_combout ;
wire \refresh_counter[11]~q ;
wire \Add0~23 ;
wire \Add0~24_combout ;
wire \refresh_counter~1_combout ;
wire \refresh_counter[12]~q ;
wire \Add0~25 ;
wire \Add0~26_combout ;
wire \refresh_counter~0_combout ;
wire \refresh_counter[13]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \i_next.000~0_combout ;
wire \i_next.000~q ;
wire \Selector7~0_combout ;
wire \i_state.000~q ;
wire \Selector8~0_combout ;
wire \i_state.001~q ;
wire \Selector16~0_combout ;
wire \Selector6~0_combout ;
wire \i_refs[0]~q ;
wire \Selector5~0_combout ;
wire \i_refs[1]~q ;
wire \Selector4~0_combout ;
wire \Selector4~1_combout ;
wire \i_refs[2]~q ;
wire \Selector18~1_combout ;
wire \Selector16~1_combout ;
wire \i_next.010~q ;
wire \Selector18~0_combout ;
wire \Selector18~2_combout ;
wire \i_next.111~q ;
wire \Selector15~1_combout ;
wire \Selector13~0_combout ;
wire \Selector15~0_combout ;
wire \Selector15~2_combout ;
wire \i_count[0]~q ;
wire \Selector14~0_combout ;
wire \Selector14~1_combout ;
wire \i_count[1]~q ;
wire \Selector12~0_combout ;
wire \i_state.111~q ;
wire \Selector13~1_combout ;
wire \Selector13~2_combout ;
wire \i_count[2]~q ;
wire \Selector9~1_combout ;
wire \i_state.010~q ;
wire \Selector10~2_combout ;
wire \Selector10~3_combout ;
wire \i_state.011~q ;
wire \Selector9~0_combout ;
wire \WideOr6~0_combout ;
wire \Selector17~0_combout ;
wire \i_next.101~q ;
wire \i_state.101~0_combout ;
wire \i_state.101~q ;
wire \init_done~0_combout ;
wire \init_done~q ;
wire \active_rnw~q ;
wire \active_addr[9]~q ;
wire \pending~0_combout ;
wire \active_addr[23]~q ;
wire \pending~1_combout ;
wire \active_addr[11]~q ;
wire \active_addr[12]~q ;
wire \pending~2_combout ;
wire \active_addr[13]~q ;
wire \active_addr[14]~q ;
wire \pending~3_combout ;
wire \pending~4_combout ;
wire \active_addr[15]~q ;
wire \active_addr[16]~q ;
wire \pending~5_combout ;
wire \active_addr[17]~q ;
wire \active_addr[18]~q ;
wire \pending~6_combout ;
wire \active_addr[19]~q ;
wire \active_addr[20]~q ;
wire \pending~7_combout ;
wire \active_addr[21]~q ;
wire \active_addr[22]~q ;
wire \pending~8_combout ;
wire \pending~9_combout ;
wire \Selector30~2_combout ;
wire \active_cs_n~0_combout ;
wire \active_cs_n~1_combout ;
wire \active_cs_n~q ;
wire \Selector41~0_combout ;
wire \Selector32~1_combout ;
wire \Selector32~0_combout ;
wire \Selector32~2_combout ;
wire \m_state.100000000~q ;
wire \pending~10_combout ;
wire \m_next~19_combout ;
wire \Selector29~0_combout ;
wire \Selector29~1_combout ;
wire \m_state.000100000~q ;
wire \Selector39~2_combout ;
wire \Selector39~3_combout ;
wire \Selector39~4_combout ;
wire \Selector39~5_combout ;
wire \Selector39~6_combout ;
wire \m_count[0]~q ;
wire \m_count~0_combout ;
wire \Selector38~0_combout ;
wire \Selector38~1_combout ;
wire \Selector38~2_combout ;
wire \Selector38~3_combout ;
wire \Selector38~4_combout ;
wire \Selector38~5_combout ;
wire \m_count[1]~q ;
wire \LessThan1~0_combout ;
wire \Selector27~0_combout ;
wire \Selector35~0_combout ;
wire \Selector25~4_combout ;
wire \Selector25~5_combout ;
wire \m_state.000000010~q ;
wire \Selector34~1_combout ;
wire \Selector34~2_combout ;
wire \Selector34~3_combout ;
wire \m_next.000010000~q ;
wire \Selector27~1_combout ;
wire \Selector28~0_combout ;
wire \Selector27~3_combout ;
wire \Selector27~4_combout ;
wire \Selector27~5_combout ;
wire \WideOr8~0_combout ;
wire \Selector27~6_combout ;
wire \m_state.000010000~q ;
wire \Selector39~7_combout ;
wire \Selector37~0_combout ;
wire \Selector37~1_combout ;
wire \Selector37~2_combout ;
wire \Selector37~3_combout ;
wire \m_count[2]~q ;
wire \Selector30~3_combout ;
wire \m_state.001000000~q ;
wire \Selector36~0_combout ;
wire \Selector36~1_combout ;
wire \Selector36~2_combout ;
wire \m_next.010000000~q ;
wire \Selector31~0_combout ;
wire \m_state.010000000~q ;
wire \Selector34~0_combout ;
wire \m_next.000001000~q ;
wire \Selector27~2_combout ;
wire \m_state.000001000~q ;
wire \WideOr9~0_combout ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \Selector26~2_combout ;
wire \m_state.000000100~q ;
wire \Selector33~0_combout ;
wire \m_addr[1]~3_combout ;
wire \Selector33~1_combout ;
wire \Selector33~2_combout ;
wire \Selector33~3_combout ;
wire \Selector33~4_combout ;
wire \m_next.000000001~q ;
wire \Selector24~0_combout ;
wire \Selector24~1_combout ;
wire \m_state.000000001~q ;
wire \Selector23~0_combout ;
wire \ack_refresh_request~q ;
wire \refresh_request~0_combout ;
wire \refresh_request~q ;
wire \active_rnw~0_combout ;
wire \active_rnw~1_combout ;
wire \active_rnw~2_combout ;
wire \active_addr[10]~q ;
wire \Selector41~1_combout ;
wire \Selector41~2_combout ;
wire \f_pop~q ;
wire \m_addr[1]~2_combout ;
wire \active_addr[0]~q ;
wire \i_addr[12]~q ;
wire \Selector97~0_combout ;
wire \Selector97~1_combout ;
wire \m_addr[1]~4_combout ;
wire \active_addr[1]~q ;
wire \Selector96~0_combout ;
wire \Selector96~1_combout ;
wire \active_addr[2]~q ;
wire \Selector95~0_combout ;
wire \Selector95~1_combout ;
wire \active_addr[3]~q ;
wire \Selector94~0_combout ;
wire \Selector94~1_combout ;
wire \active_addr[4]~q ;
wire \Selector93~0_combout ;
wire \Selector93~1_combout ;
wire \active_addr[5]~q ;
wire \f_select~combout ;
wire \Selector92~0_combout ;
wire \Selector92~1_combout ;
wire \active_addr[6]~q ;
wire \Selector91~0_combout ;
wire \Selector91~1_combout ;
wire \active_addr[7]~q ;
wire \Selector90~0_combout ;
wire \Selector90~1_combout ;
wire \active_addr[8]~q ;
wire \Selector89~0_combout ;
wire \Selector89~1_combout ;
wire \always5~0_combout ;
wire \Selector88~2_combout ;
wire \Selector88~3_combout ;
wire \Selector87~2_combout ;
wire \Selector87~3_combout ;
wire \Selector86~2_combout ;
wire \Selector86~3_combout ;
wire \Selector85~2_combout ;
wire \Selector85~3_combout ;
wire \Selector99~0_combout ;
wire \WideOr16~0_combout ;
wire \Selector98~0_combout ;
wire \Selector2~0_combout ;
wire \i_cmd[1]~q ;
wire \Selector21~0_combout ;
wire \Selector21~1_combout ;
wire \Selector0~0_combout ;
wire \i_cmd[3]~q ;
wire \Selector19~0_combout ;
wire \Selector19~1_combout ;
wire \Selector19~2_combout ;
wire \Selector19~3_combout ;
wire \active_dqm[0]~q ;
wire \Selector117~0_combout ;
wire \active_dqm[1]~q ;
wire \Selector116~0_combout ;
wire \Selector1~0_combout ;
wire \i_cmd[2]~q ;
wire \Selector20~0_combout ;
wire \Selector3~0_combout ;
wire \i_cmd[0]~q ;
wire \Selector22~0_combout ;
wire \Selector22~1_combout ;
wire \active_data[0]~q ;
wire \Selector115~0_combout ;
wire \m_data[1]~0_combout ;
wire \Selector115~1_combout ;
wire \active_data[1]~q ;
wire \Selector114~0_combout ;
wire \Selector114~1_combout ;
wire \active_data[2]~q ;
wire \Selector113~0_combout ;
wire \Selector113~1_combout ;
wire \active_data[3]~q ;
wire \Selector112~0_combout ;
wire \Selector112~1_combout ;
wire \active_data[4]~q ;
wire \Selector111~0_combout ;
wire \Selector111~1_combout ;
wire \active_data[5]~q ;
wire \Selector110~0_combout ;
wire \Selector110~1_combout ;
wire \active_data[6]~q ;
wire \Selector109~0_combout ;
wire \Selector109~1_combout ;
wire \active_data[7]~q ;
wire \Selector108~0_combout ;
wire \Selector108~1_combout ;
wire \active_data[8]~q ;
wire \Selector107~0_combout ;
wire \Selector107~1_combout ;
wire \active_data[9]~q ;
wire \Selector106~0_combout ;
wire \Selector106~1_combout ;
wire \active_data[10]~q ;
wire \Selector105~0_combout ;
wire \Selector105~1_combout ;
wire \active_data[11]~q ;
wire \Selector104~0_combout ;
wire \Selector104~1_combout ;
wire \active_data[12]~q ;
wire \Selector103~0_combout ;
wire \Selector103~1_combout ;
wire \active_data[13]~q ;
wire \Selector102~0_combout ;
wire \Selector102~1_combout ;
wire \active_data[14]~q ;
wire \Selector101~0_combout ;
wire \Selector101~1_combout ;
wire \active_data[15]~q ;
wire \Selector100~0_combout ;
wire \Selector100~1_combout ;
wire \Equal4~0_combout ;
wire \rd_valid[0]~q ;
wire \rd_valid[1]~q ;
wire \rd_valid[2]~q ;


niosII_niosII_sdram_input_efifo_module the_niosII_sdram_input_efifo_module(
	.clk(wire_pll7_clk_0),
	.reset_n(r_sync_rst),
	.f_pop(\f_pop~q ),
	.entries_1(entries_1),
	.entries_0(entries_0),
	.Equal1(\the_niosII_sdram_input_efifo_module|Equal1~0_combout ),
	.rd_data_27(\the_niosII_sdram_input_efifo_module|rd_data[27]~0_combout ),
	.rd_data_42(\the_niosII_sdram_input_efifo_module|rd_data[42]~1_combout ),
	.rd_data_41(\the_niosII_sdram_input_efifo_module|rd_data[41]~2_combout ),
	.rd_data_28(\the_niosII_sdram_input_efifo_module|rd_data[28]~3_combout ),
	.rd_data_30(\the_niosII_sdram_input_efifo_module|rd_data[30]~4_combout ),
	.rd_data_29(\the_niosII_sdram_input_efifo_module|rd_data[29]~5_combout ),
	.rd_data_32(\the_niosII_sdram_input_efifo_module|rd_data[32]~6_combout ),
	.rd_data_31(\the_niosII_sdram_input_efifo_module|rd_data[31]~7_combout ),
	.rd_data_34(\the_niosII_sdram_input_efifo_module|rd_data[34]~8_combout ),
	.rd_data_33(\the_niosII_sdram_input_efifo_module|rd_data[33]~9_combout ),
	.rd_data_36(\the_niosII_sdram_input_efifo_module|rd_data[36]~10_combout ),
	.rd_data_35(\the_niosII_sdram_input_efifo_module|rd_data[35]~11_combout ),
	.rd_data_38(\the_niosII_sdram_input_efifo_module|rd_data[38]~12_combout ),
	.rd_data_37(\the_niosII_sdram_input_efifo_module|rd_data[37]~13_combout ),
	.rd_data_40(\the_niosII_sdram_input_efifo_module|rd_data[40]~14_combout ),
	.rd_data_39(\the_niosII_sdram_input_efifo_module|rd_data[39]~15_combout ),
	.Selector41(\Selector41~0_combout ),
	.rd_data_18(\the_niosII_sdram_input_efifo_module|rd_data[18]~16_combout ),
	.rd_data_19(\the_niosII_sdram_input_efifo_module|rd_data[19]~17_combout ),
	.rd_data_20(\the_niosII_sdram_input_efifo_module|rd_data[20]~18_combout ),
	.rd_data_21(\the_niosII_sdram_input_efifo_module|rd_data[21]~19_combout ),
	.rd_data_22(\the_niosII_sdram_input_efifo_module|rd_data[22]~20_combout ),
	.rd_data_23(\the_niosII_sdram_input_efifo_module|rd_data[23]~21_combout ),
	.rd_data_24(\the_niosII_sdram_input_efifo_module|rd_data[24]~22_combout ),
	.rd_data_25(\the_niosII_sdram_input_efifo_module|rd_data[25]~23_combout ),
	.rd_data_26(\the_niosII_sdram_input_efifo_module|rd_data[26]~24_combout ),
	.rd_data_16(\the_niosII_sdram_input_efifo_module|rd_data[16]~25_combout ),
	.rd_data_17(\the_niosII_sdram_input_efifo_module|rd_data[17]~26_combout ),
	.saved_grant_0(saved_grant_0),
	.WideOr0(WideOr0),
	.Equal0(Equal0),
	.Equal11(Equal1),
	.WideOr1(WideOr1),
	.m0_write(m0_write),
	.mem_used_7(mem_used_7),
	.src_data_66(src_data_66),
	.out_data_28(out_data_28),
	.src_valid(src_valid),
	.src12_valid(src12_valid),
	.m0_write1(m0_write1),
	.out_data_42(out_data_42),
	.out_data_29(out_data_29),
	.out_data_31(out_data_31),
	.out_data_30(out_data_30),
	.out_data_33(out_data_33),
	.out_data_32(out_data_32),
	.out_data_35(out_data_35),
	.out_data_34(out_data_34),
	.out_data_37(out_data_37),
	.out_data_36(out_data_36),
	.out_data_39(out_data_39),
	.out_data_38(out_data_38),
	.out_data_41(out_data_41),
	.out_data_40(out_data_40),
	.out_data_19(out_data_19),
	.out_data_20(out_data_20),
	.out_data_21(out_data_21),
	.out_data_22(out_data_22),
	.out_data_23(out_data_23),
	.out_data_24(out_data_24),
	.out_data_25(out_data_25),
	.out_data_26(out_data_26),
	.out_data_27(out_data_27),
	.comb(\comb~1_combout ),
	.comb1(\comb~3_combout ),
	.rd_data_0(\the_niosII_sdram_input_efifo_module|rd_data[0]~27_combout ),
	.rd_data_1(\the_niosII_sdram_input_efifo_module|rd_data[1]~28_combout ),
	.rd_data_2(\the_niosII_sdram_input_efifo_module|rd_data[2]~29_combout ),
	.rd_data_3(\the_niosII_sdram_input_efifo_module|rd_data[3]~30_combout ),
	.rd_data_4(\the_niosII_sdram_input_efifo_module|rd_data[4]~31_combout ),
	.rd_data_5(\the_niosII_sdram_input_efifo_module|rd_data[5]~32_combout ),
	.rd_data_6(\the_niosII_sdram_input_efifo_module|rd_data[6]~33_combout ),
	.rd_data_7(\the_niosII_sdram_input_efifo_module|rd_data[7]~34_combout ),
	.rd_data_8(\the_niosII_sdram_input_efifo_module|rd_data[8]~35_combout ),
	.rd_data_9(\the_niosII_sdram_input_efifo_module|rd_data[9]~36_combout ),
	.rd_data_10(\the_niosII_sdram_input_efifo_module|rd_data[10]~37_combout ),
	.rd_data_11(\the_niosII_sdram_input_efifo_module|rd_data[11]~38_combout ),
	.rd_data_12(\the_niosII_sdram_input_efifo_module|rd_data[12]~39_combout ),
	.rd_data_13(\the_niosII_sdram_input_efifo_module|rd_data[13]~40_combout ),
	.rd_data_14(\the_niosII_sdram_input_efifo_module|rd_data[14]~41_combout ),
	.rd_data_15(\the_niosII_sdram_input_efifo_module|rd_data[15]~42_combout ),
	.out_data_0(out_data_0),
	.out_data_1(out_data_1),
	.out_data_2(out_data_2),
	.out_data_3(out_data_3),
	.out_data_4(out_data_4),
	.out_data_5(out_data_5),
	.out_data_6(out_data_6),
	.out_data_7(out_data_7),
	.out_data_8(out_data_8),
	.out_data_9(out_data_9),
	.out_data_10(out_data_10),
	.out_data_11(out_data_11),
	.out_data_12(out_data_12),
	.out_data_13(out_data_13),
	.out_data_14(out_data_14),
	.out_data_15(out_data_15),
	.f_select(\f_select~combout ));

cycloneive_lcell_comb \comb~0 (
	.dataa(saved_grant_1),
	.datab(d_byteenable_0),
	.datac(saved_grant_0),
	.datad(use_reg),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hFEFF;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~1 (
	.dataa(\comb~0_combout ),
	.datab(use_reg),
	.datac(byteen_reg_0),
	.datad(m0_write1),
	.cin(gnd),
	.combout(\comb~1_combout ),
	.cout());
defparam \comb~1 .lut_mask = 16'h7FFF;
defparam \comb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~2 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_1),
	.datad(use_reg),
	.cin(gnd),
	.combout(\comb~2_combout ),
	.cout());
defparam \comb~2 .lut_mask = 16'hFEFF;
defparam \comb~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~3 (
	.dataa(\comb~2_combout ),
	.datab(use_reg),
	.datac(byteen_reg_1),
	.datad(m0_write1),
	.cin(gnd),
	.combout(\comb~3_combout ),
	.cout());
defparam \comb~3 .lut_mask = 16'h7FFF;
defparam \comb~3 .sum_lutc_input = "datac";

dffeas \m_addr[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector97~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_0),
	.prn(vcc));
defparam \m_addr[0] .is_wysiwyg = "true";
defparam \m_addr[0] .power_up = "low";

dffeas \m_addr[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector96~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_1),
	.prn(vcc));
defparam \m_addr[1] .is_wysiwyg = "true";
defparam \m_addr[1] .power_up = "low";

dffeas \m_addr[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector95~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_2),
	.prn(vcc));
defparam \m_addr[2] .is_wysiwyg = "true";
defparam \m_addr[2] .power_up = "low";

dffeas \m_addr[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector94~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_3),
	.prn(vcc));
defparam \m_addr[3] .is_wysiwyg = "true";
defparam \m_addr[3] .power_up = "low";

dffeas \m_addr[4] (
	.clk(wire_pll7_clk_0),
	.d(\Selector93~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_4),
	.prn(vcc));
defparam \m_addr[4] .is_wysiwyg = "true";
defparam \m_addr[4] .power_up = "low";

dffeas \m_addr[5] (
	.clk(wire_pll7_clk_0),
	.d(\Selector92~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_5),
	.prn(vcc));
defparam \m_addr[5] .is_wysiwyg = "true";
defparam \m_addr[5] .power_up = "low";

dffeas \m_addr[6] (
	.clk(wire_pll7_clk_0),
	.d(\Selector91~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_6),
	.prn(vcc));
defparam \m_addr[6] .is_wysiwyg = "true";
defparam \m_addr[6] .power_up = "low";

dffeas \m_addr[7] (
	.clk(wire_pll7_clk_0),
	.d(\Selector90~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_7),
	.prn(vcc));
defparam \m_addr[7] .is_wysiwyg = "true";
defparam \m_addr[7] .power_up = "low";

dffeas \m_addr[8] (
	.clk(wire_pll7_clk_0),
	.d(\Selector89~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_8),
	.prn(vcc));
defparam \m_addr[8] .is_wysiwyg = "true";
defparam \m_addr[8] .power_up = "low";

dffeas oe(
	.clk(wire_pll7_clk_0),
	.d(\always5~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\m_state.000010000~q ),
	.sload(gnd),
	.ena(vcc),
	.q(oe1),
	.prn(vcc));
defparam oe.is_wysiwyg = "true";
defparam oe.power_up = "low";

dffeas \m_addr[9] (
	.clk(wire_pll7_clk_0),
	.d(\Selector88~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_9),
	.prn(vcc));
defparam \m_addr[9] .is_wysiwyg = "true";
defparam \m_addr[9] .power_up = "low";

dffeas \m_addr[10] (
	.clk(wire_pll7_clk_0),
	.d(\Selector87~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_10),
	.prn(vcc));
defparam \m_addr[10] .is_wysiwyg = "true";
defparam \m_addr[10] .power_up = "low";

dffeas \m_addr[11] (
	.clk(wire_pll7_clk_0),
	.d(\Selector86~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_11),
	.prn(vcc));
defparam \m_addr[11] .is_wysiwyg = "true";
defparam \m_addr[11] .power_up = "low";

dffeas \m_addr[12] (
	.clk(wire_pll7_clk_0),
	.d(\Selector85~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[1]~4_combout ),
	.q(m_addr_12),
	.prn(vcc));
defparam \m_addr[12] .is_wysiwyg = "true";
defparam \m_addr[12] .power_up = "low";

dffeas \m_bank[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector99~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_bank_0),
	.prn(vcc));
defparam \m_bank[0] .is_wysiwyg = "true";
defparam \m_bank[0] .power_up = "low";

dffeas \m_bank[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector98~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_bank_1),
	.prn(vcc));
defparam \m_bank[1] .is_wysiwyg = "true";
defparam \m_bank[1] .power_up = "low";

dffeas \m_cmd[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector21~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_1),
	.prn(vcc));
defparam \m_cmd[1] .is_wysiwyg = "true";
defparam \m_cmd[1] .power_up = "low";

dffeas \m_cmd[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector19~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_3),
	.prn(vcc));
defparam \m_cmd[3] .is_wysiwyg = "true";
defparam \m_cmd[3] .power_up = "low";

dffeas \m_dqm[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector117~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_0),
	.prn(vcc));
defparam \m_dqm[0] .is_wysiwyg = "true";
defparam \m_dqm[0] .power_up = "low";

dffeas \m_dqm[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector116~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_1),
	.prn(vcc));
defparam \m_dqm[1] .is_wysiwyg = "true";
defparam \m_dqm[1] .power_up = "low";

dffeas \m_cmd[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_2),
	.prn(vcc));
defparam \m_cmd[2] .is_wysiwyg = "true";
defparam \m_cmd[2] .power_up = "low";

dffeas \m_cmd[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector22~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_0),
	.prn(vcc));
defparam \m_cmd[0] .is_wysiwyg = "true";
defparam \m_cmd[0] .power_up = "low";

dffeas \m_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector115~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_0),
	.prn(vcc));
defparam \m_data[0] .is_wysiwyg = "true";
defparam \m_data[0] .power_up = "low";

dffeas \m_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector114~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_1),
	.prn(vcc));
defparam \m_data[1] .is_wysiwyg = "true";
defparam \m_data[1] .power_up = "low";

dffeas \m_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector113~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_2),
	.prn(vcc));
defparam \m_data[2] .is_wysiwyg = "true";
defparam \m_data[2] .power_up = "low";

dffeas \m_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector112~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_3),
	.prn(vcc));
defparam \m_data[3] .is_wysiwyg = "true";
defparam \m_data[3] .power_up = "low";

dffeas \m_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\Selector111~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_4),
	.prn(vcc));
defparam \m_data[4] .is_wysiwyg = "true";
defparam \m_data[4] .power_up = "low";

dffeas \m_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\Selector110~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_5),
	.prn(vcc));
defparam \m_data[5] .is_wysiwyg = "true";
defparam \m_data[5] .power_up = "low";

dffeas \m_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\Selector109~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_6),
	.prn(vcc));
defparam \m_data[6] .is_wysiwyg = "true";
defparam \m_data[6] .power_up = "low";

dffeas \m_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\Selector108~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_7),
	.prn(vcc));
defparam \m_data[7] .is_wysiwyg = "true";
defparam \m_data[7] .power_up = "low";

dffeas \m_data[8] (
	.clk(wire_pll7_clk_0),
	.d(\Selector107~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_8),
	.prn(vcc));
defparam \m_data[8] .is_wysiwyg = "true";
defparam \m_data[8] .power_up = "low";

dffeas \m_data[9] (
	.clk(wire_pll7_clk_0),
	.d(\Selector106~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_9),
	.prn(vcc));
defparam \m_data[9] .is_wysiwyg = "true";
defparam \m_data[9] .power_up = "low";

dffeas \m_data[10] (
	.clk(wire_pll7_clk_0),
	.d(\Selector105~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_10),
	.prn(vcc));
defparam \m_data[10] .is_wysiwyg = "true";
defparam \m_data[10] .power_up = "low";

dffeas \m_data[11] (
	.clk(wire_pll7_clk_0),
	.d(\Selector104~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_11),
	.prn(vcc));
defparam \m_data[11] .is_wysiwyg = "true";
defparam \m_data[11] .power_up = "low";

dffeas \m_data[12] (
	.clk(wire_pll7_clk_0),
	.d(\Selector103~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_12),
	.prn(vcc));
defparam \m_data[12] .is_wysiwyg = "true";
defparam \m_data[12] .power_up = "low";

dffeas \m_data[13] (
	.clk(wire_pll7_clk_0),
	.d(\Selector102~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_13),
	.prn(vcc));
defparam \m_data[13] .is_wysiwyg = "true";
defparam \m_data[13] .power_up = "low";

dffeas \m_data[14] (
	.clk(wire_pll7_clk_0),
	.d(\Selector101~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_14),
	.prn(vcc));
defparam \m_data[14] .is_wysiwyg = "true";
defparam \m_data[14] .power_up = "low";

dffeas \m_data[15] (
	.clk(wire_pll7_clk_0),
	.d(\Selector100~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_15),
	.prn(vcc));
defparam \m_data[15] .is_wysiwyg = "true";
defparam \m_data[15] .power_up = "low";

dffeas za_valid(
	.clk(wire_pll7_clk_0),
	.d(\rd_valid[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_valid1),
	.prn(vcc));
defparam za_valid.is_wysiwyg = "true";
defparam za_valid.power_up = "low";

dffeas \za_data[0] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_0),
	.prn(vcc));
defparam \za_data[0] .is_wysiwyg = "true";
defparam \za_data[0] .power_up = "low";

dffeas \za_data[1] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_1),
	.prn(vcc));
defparam \za_data[1] .is_wysiwyg = "true";
defparam \za_data[1] .power_up = "low";

dffeas \za_data[2] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_2),
	.prn(vcc));
defparam \za_data[2] .is_wysiwyg = "true";
defparam \za_data[2] .power_up = "low";

dffeas \za_data[3] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_3),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_3),
	.prn(vcc));
defparam \za_data[3] .is_wysiwyg = "true";
defparam \za_data[3] .power_up = "low";

dffeas \za_data[4] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_4),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_4),
	.prn(vcc));
defparam \za_data[4] .is_wysiwyg = "true";
defparam \za_data[4] .power_up = "low";

dffeas \za_data[11] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_11),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_11),
	.prn(vcc));
defparam \za_data[11] .is_wysiwyg = "true";
defparam \za_data[11] .power_up = "low";

dffeas \za_data[13] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_13),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_13),
	.prn(vcc));
defparam \za_data[13] .is_wysiwyg = "true";
defparam \za_data[13] .power_up = "low";

dffeas \za_data[12] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_12),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_12),
	.prn(vcc));
defparam \za_data[12] .is_wysiwyg = "true";
defparam \za_data[12] .power_up = "low";

dffeas \za_data[5] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_5),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_5),
	.prn(vcc));
defparam \za_data[5] .is_wysiwyg = "true";
defparam \za_data[5] .power_up = "low";

dffeas \za_data[14] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_14),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_14),
	.prn(vcc));
defparam \za_data[14] .is_wysiwyg = "true";
defparam \za_data[14] .power_up = "low";

dffeas \za_data[15] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_15),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_15),
	.prn(vcc));
defparam \za_data[15] .is_wysiwyg = "true";
defparam \za_data[15] .power_up = "low";

dffeas \za_data[10] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_10),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_10),
	.prn(vcc));
defparam \za_data[10] .is_wysiwyg = "true";
defparam \za_data[10] .power_up = "low";

dffeas \za_data[9] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_9),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_9),
	.prn(vcc));
defparam \za_data[9] .is_wysiwyg = "true";
defparam \za_data[9] .power_up = "low";

dffeas \za_data[8] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_8),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_8),
	.prn(vcc));
defparam \za_data[8] .is_wysiwyg = "true";
defparam \za_data[8] .power_up = "low";

dffeas \za_data[7] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_7),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_7),
	.prn(vcc));
defparam \za_data[7] .is_wysiwyg = "true";
defparam \za_data[7] .power_up = "low";

dffeas \za_data[6] (
	.clk(wire_pll7_clk_0),
	.d(sdram_dq_6),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_6),
	.prn(vcc));
defparam \za_data[6] .is_wysiwyg = "true";
defparam \za_data[6] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(\refresh_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh_counter~8 (
	.dataa(\Add0~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~8_combout ),
	.cout());
defparam \refresh_counter~8 .lut_mask = 16'hAAFF;
defparam \refresh_counter~8 .sum_lutc_input = "datac";

dffeas \refresh_counter[0] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[0]~q ),
	.prn(vcc));
defparam \refresh_counter[0] .is_wysiwyg = "true";
defparam \refresh_counter[0] .power_up = "low";

cycloneive_lcell_comb \Add0~2 (
	.dataa(\refresh_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

dffeas \refresh_counter[1] (
	.clk(wire_pll7_clk_0),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[1]~q ),
	.prn(vcc));
defparam \refresh_counter[1] .is_wysiwyg = "true";
defparam \refresh_counter[1] .power_up = "low";

cycloneive_lcell_comb \Add0~4 (
	.dataa(\refresh_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~7 (
	.dataa(\Add0~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~7_combout ),
	.cout());
defparam \refresh_counter~7 .lut_mask = 16'hAAFF;
defparam \refresh_counter~7 .sum_lutc_input = "datac";

dffeas \refresh_counter[2] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[2]~q ),
	.prn(vcc));
defparam \refresh_counter[2] .is_wysiwyg = "true";
defparam \refresh_counter[2] .power_up = "low";

cycloneive_lcell_comb \Add0~6 (
	.dataa(\refresh_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

dffeas \refresh_counter[3] (
	.clk(wire_pll7_clk_0),
	.d(\Add0~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[3]~q ),
	.prn(vcc));
defparam \refresh_counter[3] .is_wysiwyg = "true";
defparam \refresh_counter[3] .power_up = "low";

cycloneive_lcell_comb \Add0~8 (
	.dataa(\refresh_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5A5F;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter[4]~13 (
	.dataa(\Add0~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\refresh_counter[4]~13_combout ),
	.cout());
defparam \refresh_counter[4]~13 .lut_mask = 16'h5555;
defparam \refresh_counter[4]~13 .sum_lutc_input = "datac";

dffeas \refresh_counter[4] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter[4]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[4]~q ),
	.prn(vcc));
defparam \refresh_counter[4] .is_wysiwyg = "true";
defparam \refresh_counter[4] .power_up = "low";

cycloneive_lcell_comb \Add0~10 (
	.dataa(\refresh_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~6 (
	.dataa(\Add0~10_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~6_combout ),
	.cout());
defparam \refresh_counter~6 .lut_mask = 16'hAAFF;
defparam \refresh_counter~6 .sum_lutc_input = "datac";

dffeas \refresh_counter[5] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[5]~q ),
	.prn(vcc));
defparam \refresh_counter[5] .is_wysiwyg = "true";
defparam \refresh_counter[5] .power_up = "low";

cycloneive_lcell_comb \Add0~12 (
	.dataa(\refresh_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5AAF;
defparam \Add0~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~5 (
	.dataa(\Add0~12_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~5_combout ),
	.cout());
defparam \refresh_counter~5 .lut_mask = 16'hAAFF;
defparam \refresh_counter~5 .sum_lutc_input = "datac";

dffeas \refresh_counter[6] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[6]~q ),
	.prn(vcc));
defparam \refresh_counter[6] .is_wysiwyg = "true";
defparam \refresh_counter[6] .power_up = "low";

cycloneive_lcell_comb \Add0~14 (
	.dataa(\refresh_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~4 (
	.dataa(\Add0~14_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~4_combout ),
	.cout());
defparam \refresh_counter~4 .lut_mask = 16'hAAFF;
defparam \refresh_counter~4 .sum_lutc_input = "datac";

dffeas \refresh_counter[7] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[7]~q ),
	.prn(vcc));
defparam \refresh_counter[7] .is_wysiwyg = "true";
defparam \refresh_counter[7] .power_up = "low";

cycloneive_lcell_comb \Add0~16 (
	.dataa(\refresh_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
defparam \Add0~16 .lut_mask = 16'h5A5F;
defparam \Add0~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~3 (
	.dataa(\Add0~16_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~3_combout ),
	.cout());
defparam \refresh_counter~3 .lut_mask = 16'hFF55;
defparam \refresh_counter~3 .sum_lutc_input = "datac";

dffeas \refresh_counter[8] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[8]~q ),
	.prn(vcc));
defparam \refresh_counter[8] .is_wysiwyg = "true";
defparam \refresh_counter[8] .power_up = "low";

cycloneive_lcell_comb \Add0~18 (
	.dataa(\refresh_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
defparam \Add0~18 .lut_mask = 16'h5AAF;
defparam \Add0~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter[9]~11 (
	.dataa(\Add0~18_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\refresh_counter[9]~11_combout ),
	.cout());
defparam \refresh_counter[9]~11 .lut_mask = 16'h5555;
defparam \refresh_counter[9]~11 .sum_lutc_input = "datac";

dffeas \refresh_counter[9] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter[9]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[9]~q ),
	.prn(vcc));
defparam \refresh_counter[9] .is_wysiwyg = "true";
defparam \refresh_counter[9] .power_up = "low";

cycloneive_lcell_comb \Add0~20 (
	.dataa(\refresh_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
defparam \Add0~20 .lut_mask = 16'h5A5F;
defparam \Add0~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter[10]~10 (
	.dataa(\Add0~20_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\refresh_counter[10]~10_combout ),
	.cout());
defparam \refresh_counter[10]~10 .lut_mask = 16'h5555;
defparam \refresh_counter[10]~10 .sum_lutc_input = "datac";

dffeas \refresh_counter[10] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter[10]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[10]~q ),
	.prn(vcc));
defparam \refresh_counter[10] .is_wysiwyg = "true";
defparam \refresh_counter[10] .power_up = "low";

cycloneive_lcell_comb \Add0~22 (
	.dataa(\refresh_counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
defparam \Add0~22 .lut_mask = 16'h5A5F;
defparam \Add0~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~2 (
	.dataa(\Add0~22_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~2_combout ),
	.cout());
defparam \refresh_counter~2 .lut_mask = 16'hAAFF;
defparam \refresh_counter~2 .sum_lutc_input = "datac";

dffeas \refresh_counter[11] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[11]~q ),
	.prn(vcc));
defparam \refresh_counter[11] .is_wysiwyg = "true";
defparam \refresh_counter[11] .power_up = "low";

cycloneive_lcell_comb \Add0~24 (
	.dataa(\refresh_counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
defparam \Add0~24 .lut_mask = 16'h5AAF;
defparam \Add0~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~1 (
	.dataa(\Add0~24_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~1_combout ),
	.cout());
defparam \refresh_counter~1 .lut_mask = 16'hAAFF;
defparam \refresh_counter~1 .sum_lutc_input = "datac";

dffeas \refresh_counter[12] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[12]~q ),
	.prn(vcc));
defparam \refresh_counter[12] .is_wysiwyg = "true";
defparam \refresh_counter[12] .power_up = "low";

cycloneive_lcell_comb \Add0~26 (
	.dataa(\refresh_counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout());
defparam \Add0~26 .lut_mask = 16'h5A5A;
defparam \Add0~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~0 (
	.dataa(\Add0~26_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~0_combout ),
	.cout());
defparam \refresh_counter~0 .lut_mask = 16'hFF55;
defparam \refresh_counter~0 .sum_lutc_input = "datac";

dffeas \refresh_counter[13] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[13]~q ),
	.prn(vcc));
defparam \refresh_counter[13] .is_wysiwyg = "true";
defparam \refresh_counter[13] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\refresh_counter[13]~q ),
	.datab(\refresh_counter[10]~q ),
	.datac(\refresh_counter[12]~q ),
	.datad(\refresh_counter[11]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\refresh_counter[9]~q ),
	.datab(\refresh_counter[8]~q ),
	.datac(\refresh_counter[7]~q ),
	.datad(\refresh_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\refresh_counter[4]~q ),
	.datab(\refresh_counter[5]~q ),
	.datac(\refresh_counter[3]~q ),
	.datad(\refresh_counter[2]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hBFFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\refresh_counter[1]~q ),
	.datad(\refresh_counter[0]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'h0FFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'hFFFE;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_next.000~0 (
	.dataa(\i_next.000~q ),
	.datab(\i_state.000~q ),
	.datac(\i_state.101~q ),
	.datad(\i_state.011~q ),
	.cin(gnd),
	.combout(\i_next.000~0_combout ),
	.cout());
defparam \i_next.000~0 .lut_mask = 16'hEFFF;
defparam \i_next.000~0 .sum_lutc_input = "datac";

dffeas \i_next.000 (
	.clk(wire_pll7_clk_0),
	.d(\i_next.000~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.000~q ),
	.prn(vcc));
defparam \i_next.000 .is_wysiwyg = "true";
defparam \i_next.000 .power_up = "low";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(\Selector9~0_combout ),
	.datab(\i_state.000~q ),
	.datac(\Equal0~4_combout ),
	.datad(\i_next.000~q ),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hFFFD;
defparam \Selector7~0 .sum_lutc_input = "datac";

dffeas \i_state.000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.000~q ),
	.prn(vcc));
defparam \i_state.000 .is_wysiwyg = "true";
defparam \i_state.000 .power_up = "low";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(\Equal0~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hAAFF;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \i_state.001 (
	.clk(wire_pll7_clk_0),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.001~q ),
	.prn(vcc));
defparam \i_state.001 .is_wysiwyg = "true";
defparam \i_state.001 .power_up = "low";

cycloneive_lcell_comb \Selector16~0 (
	.dataa(\i_next.010~q ),
	.datab(\i_state.101~q ),
	.datac(\i_state.011~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
defparam \Selector16~0 .lut_mask = 16'hFEFF;
defparam \Selector16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(\i_state.000~q ),
	.datab(gnd),
	.datac(\i_state.010~q ),
	.datad(\i_refs[0]~q ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hAFFA;
defparam \Selector6~0 .sum_lutc_input = "datac";

dffeas \i_refs[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!r_sync_rst),
	.q(\i_refs[0]~q ),
	.prn(vcc));
defparam \i_refs[0] .is_wysiwyg = "true";
defparam \i_refs[0] .power_up = "low";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\i_state.000~q ),
	.datab(\i_state.010~q ),
	.datac(\i_refs[1]~q ),
	.datad(\i_refs[0]~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hEBBE;
defparam \Selector5~0 .sum_lutc_input = "datac";

dffeas \i_refs[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!r_sync_rst),
	.q(\i_refs[1]~q ),
	.prn(vcc));
defparam \i_refs[1] .is_wysiwyg = "true";
defparam \i_refs[1] .power_up = "low";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(\i_state.010~q ),
	.datab(\i_refs[2]~q ),
	.datac(\i_refs[1]~q ),
	.datad(\i_refs[0]~q ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hEBBE;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~1 (
	.dataa(\Selector4~0_combout ),
	.datab(\i_state.000~q ),
	.datac(\i_refs[2]~q ),
	.datad(\i_state.010~q ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hFEFF;
defparam \Selector4~1 .sum_lutc_input = "datac";

dffeas \i_refs[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!r_sync_rst),
	.q(\i_refs[2]~q ),
	.prn(vcc));
defparam \i_refs[2] .is_wysiwyg = "true";
defparam \i_refs[2] .power_up = "low";

cycloneive_lcell_comb \Selector18~1 (
	.dataa(\i_refs[0]~q ),
	.datab(gnd),
	.datac(\i_refs[2]~q ),
	.datad(\i_refs[1]~q ),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
defparam \Selector18~1 .lut_mask = 16'hAFFF;
defparam \Selector18~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector16~1 (
	.dataa(\i_state.001~q ),
	.datab(\Selector16~0_combout ),
	.datac(\i_state.010~q ),
	.datad(\Selector18~1_combout ),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
defparam \Selector16~1 .lut_mask = 16'hFEFF;
defparam \Selector16~1 .sum_lutc_input = "datac";

dffeas \i_next.010 (
	.clk(wire_pll7_clk_0),
	.d(\Selector16~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.010~q ),
	.prn(vcc));
defparam \i_next.010 .is_wysiwyg = "true";
defparam \i_next.010 .power_up = "low";

cycloneive_lcell_comb \Selector18~0 (
	.dataa(\i_next.111~q ),
	.datab(\i_state.101~q ),
	.datac(\i_state.011~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
defparam \Selector18~0 .lut_mask = 16'hFEFF;
defparam \Selector18~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector18~2 (
	.dataa(\Selector18~0_combout ),
	.datab(\i_state.010~q ),
	.datac(\Selector18~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector18~2_combout ),
	.cout());
defparam \Selector18~2 .lut_mask = 16'hFEFE;
defparam \Selector18~2 .sum_lutc_input = "datac";

dffeas \i_next.111 (
	.clk(wire_pll7_clk_0),
	.d(\Selector18~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.111~q ),
	.prn(vcc));
defparam \i_next.111 .is_wysiwyg = "true";
defparam \i_next.111 .power_up = "low";

cycloneive_lcell_comb \Selector15~1 (
	.dataa(\i_state.011~q ),
	.datab(\i_count[2]~q ),
	.datac(\i_count[1]~q ),
	.datad(\i_count[0]~q ),
	.cin(gnd),
	.combout(\Selector15~1_combout ),
	.cout());
defparam \Selector15~1 .lut_mask = 16'hEBBE;
defparam \Selector15~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector13~0 (
	.dataa(\i_state.000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\i_state.101~q ),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
defparam \Selector13~0 .lut_mask = 16'hAAFF;
defparam \Selector13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector15~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\i_state.001~q ),
	.datad(\i_state.010~q ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
defparam \Selector15~0 .lut_mask = 16'h0FFF;
defparam \Selector15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector15~2 (
	.dataa(\Selector15~1_combout ),
	.datab(\i_count[0]~q ),
	.datac(\Selector13~0_combout ),
	.datad(\Selector15~0_combout ),
	.cin(gnd),
	.combout(\Selector15~2_combout ),
	.cout());
defparam \Selector15~2 .lut_mask = 16'hEFFF;
defparam \Selector15~2 .sum_lutc_input = "datac";

dffeas \i_count[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector15~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[0]~q ),
	.prn(vcc));
defparam \i_count[0] .is_wysiwyg = "true";
defparam \i_count[0] .power_up = "low";

cycloneive_lcell_comb \Selector14~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_count[1]~q ),
	.datac(\i_count[0]~q ),
	.datad(\i_count[2]~q ),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
defparam \Selector14~0 .lut_mask = 16'hFFBE;
defparam \Selector14~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector14~1 (
	.dataa(\i_state.010~q ),
	.datab(\Selector14~0_combout ),
	.datac(\i_count[1]~q ),
	.datad(\Selector13~0_combout ),
	.cin(gnd),
	.combout(\Selector14~1_combout ),
	.cout());
defparam \Selector14~1 .lut_mask = 16'hFEFF;
defparam \Selector14~1 .sum_lutc_input = "datac";

dffeas \i_count[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector14~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[1]~q ),
	.prn(vcc));
defparam \i_count[1] .is_wysiwyg = "true";
defparam \i_count[1] .power_up = "low";

cycloneive_lcell_comb \Selector12~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_next.111~q ),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
defparam \Selector12~0 .lut_mask = 16'hEFFF;
defparam \Selector12~0 .sum_lutc_input = "datac";

dffeas \i_state.111 (
	.clk(wire_pll7_clk_0),
	.d(\Selector12~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.111~q ),
	.prn(vcc));
defparam \i_state.111 .is_wysiwyg = "true";
defparam \i_state.111 .power_up = "low";

cycloneive_lcell_comb \Selector13~1 (
	.dataa(\i_state.011~q ),
	.datab(\i_count[1]~q ),
	.datac(\i_count[0]~q ),
	.datad(\Selector13~0_combout ),
	.cin(gnd),
	.combout(\Selector13~1_combout ),
	.cout());
defparam \Selector13~1 .lut_mask = 16'hFEFF;
defparam \Selector13~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector13~2 (
	.dataa(\i_state.111~q ),
	.datab(\i_state.010~q ),
	.datac(\i_count[2]~q ),
	.datad(\Selector13~1_combout ),
	.cin(gnd),
	.combout(\Selector13~2_combout ),
	.cout());
defparam \Selector13~2 .lut_mask = 16'hFFFE;
defparam \Selector13~2 .sum_lutc_input = "datac";

dffeas \i_count[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector13~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[2]~q ),
	.prn(vcc));
defparam \i_count[2] .is_wysiwyg = "true";
defparam \i_count[2] .power_up = "low";

cycloneive_lcell_comb \Selector9~1 (
	.dataa(\i_state.011~q ),
	.datab(\i_next.010~q ),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector9~1_combout ),
	.cout());
defparam \Selector9~1 .lut_mask = 16'hEFFF;
defparam \Selector9~1 .sum_lutc_input = "datac";

dffeas \i_state.010 (
	.clk(wire_pll7_clk_0),
	.d(\Selector9~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.010~q ),
	.prn(vcc));
defparam \i_state.010 .is_wysiwyg = "true";
defparam \i_state.010 .power_up = "low";

cycloneive_lcell_comb \Selector10~2 (
	.dataa(\i_state.111~q ),
	.datab(\i_state.011~q ),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
defparam \Selector10~2 .lut_mask = 16'hFFFE;
defparam \Selector10~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector10~3 (
	.dataa(\i_state.001~q ),
	.datab(\i_state.010~q ),
	.datac(\Selector10~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector10~3_combout ),
	.cout());
defparam \Selector10~3 .lut_mask = 16'hFEFE;
defparam \Selector10~3 .sum_lutc_input = "datac";

dffeas \i_state.011 (
	.clk(wire_pll7_clk_0),
	.d(\Selector10~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.011~q ),
	.prn(vcc));
defparam \i_state.011 .is_wysiwyg = "true";
defparam \i_state.011 .power_up = "low";

cycloneive_lcell_comb \Selector9~0 (
	.dataa(\i_state.011~q ),
	.datab(gnd),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hAFFF;
defparam \Selector9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr6~0 (
	.dataa(\i_state.000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\i_state.011~q ),
	.cin(gnd),
	.combout(\WideOr6~0_combout ),
	.cout());
defparam \WideOr6~0 .lut_mask = 16'hAAFF;
defparam \WideOr6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector17~0 (
	.dataa(\i_state.111~q ),
	.datab(\i_next.101~q ),
	.datac(\i_state.101~q ),
	.datad(\WideOr6~0_combout ),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
defparam \Selector17~0 .lut_mask = 16'hFEFF;
defparam \Selector17~0 .sum_lutc_input = "datac";

dffeas \i_next.101 (
	.clk(wire_pll7_clk_0),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.101~q ),
	.prn(vcc));
defparam \i_next.101 .is_wysiwyg = "true";
defparam \i_next.101 .power_up = "low";

cycloneive_lcell_comb \i_state.101~0 (
	.dataa(\i_state.101~q ),
	.datab(\Selector9~0_combout ),
	.datac(\i_next.101~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\i_state.101~0_combout ),
	.cout());
defparam \i_state.101~0 .lut_mask = 16'hFEFE;
defparam \i_state.101~0 .sum_lutc_input = "datac";

dffeas \i_state.101 (
	.clk(wire_pll7_clk_0),
	.d(\i_state.101~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.101~q ),
	.prn(vcc));
defparam \i_state.101 .is_wysiwyg = "true";
defparam \i_state.101 .power_up = "low";

cycloneive_lcell_comb \init_done~0 (
	.dataa(\init_done~q ),
	.datab(\i_state.101~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\init_done~0_combout ),
	.cout());
defparam \init_done~0 .lut_mask = 16'hEEEE;
defparam \init_done~0 .sum_lutc_input = "datac";

dffeas init_done(
	.clk(wire_pll7_clk_0),
	.d(\init_done~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\init_done~q ),
	.prn(vcc));
defparam init_done.is_wysiwyg = "true";
defparam init_done.power_up = "low";

dffeas active_rnw(
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[42]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_rnw~q ),
	.prn(vcc));
defparam active_rnw.is_wysiwyg = "true";
defparam active_rnw.power_up = "low";

dffeas \active_addr[9] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[27]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[9]~q ),
	.prn(vcc));
defparam \active_addr[9] .is_wysiwyg = "true";
defparam \active_addr[9] .power_up = "low";

cycloneive_lcell_comb \pending~0 (
	.dataa(\active_rnw~q ),
	.datab(\active_addr[9]~q ),
	.datac(\the_niosII_sdram_input_efifo_module|rd_data[27]~0_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[42]~1_combout ),
	.cin(gnd),
	.combout(\pending~0_combout ),
	.cout());
defparam \pending~0 .lut_mask = 16'h6996;
defparam \pending~0 .sum_lutc_input = "datac";

dffeas \active_addr[23] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[41]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[23]~q ),
	.prn(vcc));
defparam \active_addr[23] .is_wysiwyg = "true";
defparam \active_addr[23] .power_up = "low";

cycloneive_lcell_comb \pending~1 (
	.dataa(\active_addr[10]~q ),
	.datab(\active_addr[23]~q ),
	.datac(\the_niosII_sdram_input_efifo_module|rd_data[41]~2_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[28]~3_combout ),
	.cin(gnd),
	.combout(\pending~1_combout ),
	.cout());
defparam \pending~1 .lut_mask = 16'h6996;
defparam \pending~1 .sum_lutc_input = "datac";

dffeas \active_addr[11] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[29]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[11]~q ),
	.prn(vcc));
defparam \active_addr[11] .is_wysiwyg = "true";
defparam \active_addr[11] .power_up = "low";

dffeas \active_addr[12] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[30]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[12]~q ),
	.prn(vcc));
defparam \active_addr[12] .is_wysiwyg = "true";
defparam \active_addr[12] .power_up = "low";

cycloneive_lcell_comb \pending~2 (
	.dataa(\active_addr[11]~q ),
	.datab(\active_addr[12]~q ),
	.datac(\the_niosII_sdram_input_efifo_module|rd_data[30]~4_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[29]~5_combout ),
	.cin(gnd),
	.combout(\pending~2_combout ),
	.cout());
defparam \pending~2 .lut_mask = 16'h6996;
defparam \pending~2 .sum_lutc_input = "datac";

dffeas \active_addr[13] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[31]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[13]~q ),
	.prn(vcc));
defparam \active_addr[13] .is_wysiwyg = "true";
defparam \active_addr[13] .power_up = "low";

dffeas \active_addr[14] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[32]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[14]~q ),
	.prn(vcc));
defparam \active_addr[14] .is_wysiwyg = "true";
defparam \active_addr[14] .power_up = "low";

cycloneive_lcell_comb \pending~3 (
	.dataa(\active_addr[13]~q ),
	.datab(\active_addr[14]~q ),
	.datac(\the_niosII_sdram_input_efifo_module|rd_data[32]~6_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[31]~7_combout ),
	.cin(gnd),
	.combout(\pending~3_combout ),
	.cout());
defparam \pending~3 .lut_mask = 16'h6996;
defparam \pending~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \pending~4 (
	.dataa(\pending~0_combout ),
	.datab(\pending~1_combout ),
	.datac(\pending~2_combout ),
	.datad(\pending~3_combout ),
	.cin(gnd),
	.combout(\pending~4_combout ),
	.cout());
defparam \pending~4 .lut_mask = 16'hFFFE;
defparam \pending~4 .sum_lutc_input = "datac";

dffeas \active_addr[15] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[33]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[15]~q ),
	.prn(vcc));
defparam \active_addr[15] .is_wysiwyg = "true";
defparam \active_addr[15] .power_up = "low";

dffeas \active_addr[16] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[34]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[16]~q ),
	.prn(vcc));
defparam \active_addr[16] .is_wysiwyg = "true";
defparam \active_addr[16] .power_up = "low";

cycloneive_lcell_comb \pending~5 (
	.dataa(\active_addr[15]~q ),
	.datab(\active_addr[16]~q ),
	.datac(\the_niosII_sdram_input_efifo_module|rd_data[34]~8_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[33]~9_combout ),
	.cin(gnd),
	.combout(\pending~5_combout ),
	.cout());
defparam \pending~5 .lut_mask = 16'h6996;
defparam \pending~5 .sum_lutc_input = "datac";

dffeas \active_addr[17] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[35]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[17]~q ),
	.prn(vcc));
defparam \active_addr[17] .is_wysiwyg = "true";
defparam \active_addr[17] .power_up = "low";

dffeas \active_addr[18] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[36]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[18]~q ),
	.prn(vcc));
defparam \active_addr[18] .is_wysiwyg = "true";
defparam \active_addr[18] .power_up = "low";

cycloneive_lcell_comb \pending~6 (
	.dataa(\active_addr[17]~q ),
	.datab(\active_addr[18]~q ),
	.datac(\the_niosII_sdram_input_efifo_module|rd_data[36]~10_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[35]~11_combout ),
	.cin(gnd),
	.combout(\pending~6_combout ),
	.cout());
defparam \pending~6 .lut_mask = 16'h6996;
defparam \pending~6 .sum_lutc_input = "datac";

dffeas \active_addr[19] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[37]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[19]~q ),
	.prn(vcc));
defparam \active_addr[19] .is_wysiwyg = "true";
defparam \active_addr[19] .power_up = "low";

dffeas \active_addr[20] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[38]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[20]~q ),
	.prn(vcc));
defparam \active_addr[20] .is_wysiwyg = "true";
defparam \active_addr[20] .power_up = "low";

cycloneive_lcell_comb \pending~7 (
	.dataa(\active_addr[19]~q ),
	.datab(\active_addr[20]~q ),
	.datac(\the_niosII_sdram_input_efifo_module|rd_data[38]~12_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[37]~13_combout ),
	.cin(gnd),
	.combout(\pending~7_combout ),
	.cout());
defparam \pending~7 .lut_mask = 16'h6996;
defparam \pending~7 .sum_lutc_input = "datac";

dffeas \active_addr[21] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[39]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[21]~q ),
	.prn(vcc));
defparam \active_addr[21] .is_wysiwyg = "true";
defparam \active_addr[21] .power_up = "low";

dffeas \active_addr[22] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[40]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[22]~q ),
	.prn(vcc));
defparam \active_addr[22] .is_wysiwyg = "true";
defparam \active_addr[22] .power_up = "low";

cycloneive_lcell_comb \pending~8 (
	.dataa(\active_addr[21]~q ),
	.datab(\active_addr[22]~q ),
	.datac(\the_niosII_sdram_input_efifo_module|rd_data[40]~14_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[39]~15_combout ),
	.cin(gnd),
	.combout(\pending~8_combout ),
	.cout());
defparam \pending~8 .lut_mask = 16'h6996;
defparam \pending~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \pending~9 (
	.dataa(\pending~5_combout ),
	.datab(\pending~6_combout ),
	.datac(\pending~7_combout ),
	.datad(\pending~8_combout ),
	.cin(gnd),
	.combout(\pending~9_combout ),
	.cout());
defparam \pending~9 .lut_mask = 16'hFFFE;
defparam \pending~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector30~2 (
	.dataa(\init_done~q ),
	.datab(\refresh_request~q ),
	.datac(gnd),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector30~2_combout ),
	.cout());
defparam \Selector30~2 .lut_mask = 16'hEEFF;
defparam \Selector30~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_cs_n~0 (
	.dataa(\m_state.000000001~q ),
	.datab(entries_1),
	.datac(entries_0),
	.datad(\init_done~q ),
	.cin(gnd),
	.combout(\active_cs_n~0_combout ),
	.cout());
defparam \active_cs_n~0 .lut_mask = 16'hBFFF;
defparam \active_cs_n~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_cs_n~1 (
	.dataa(\active_cs_n~q ),
	.datab(\Selector30~2_combout ),
	.datac(\active_cs_n~0_combout ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\active_cs_n~1_combout ),
	.cout());
defparam \active_cs_n~1 .lut_mask = 16'hFAFC;
defparam \active_cs_n~1 .sum_lutc_input = "datac";

dffeas active_cs_n(
	.clk(wire_pll7_clk_0),
	.d(\active_cs_n~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\active_cs_n~q ),
	.prn(vcc));
defparam active_cs_n.is_wysiwyg = "true";
defparam active_cs_n.power_up = "low";

cycloneive_lcell_comb \Selector41~0 (
	.dataa(\the_niosII_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(\pending~4_combout ),
	.datac(\pending~9_combout ),
	.datad(\active_cs_n~q ),
	.cin(gnd),
	.combout(\Selector41~0_combout ),
	.cout());
defparam \Selector41~0 .lut_mask = 16'hFEFF;
defparam \Selector41~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector32~1 (
	.dataa(\m_state.100000000~q ),
	.datab(\refresh_request~q ),
	.datac(\Selector41~0_combout ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector32~1_combout ),
	.cout());
defparam \Selector32~1 .lut_mask = 16'hBFFF;
defparam \Selector32~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector32~0 (
	.dataa(gnd),
	.datab(entries_1),
	.datac(entries_0),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector32~0_combout ),
	.cout());
defparam \Selector32~0 .lut_mask = 16'h3FFF;
defparam \Selector32~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector32~2 (
	.dataa(\Selector32~1_combout ),
	.datab(\m_state.100000000~q ),
	.datac(\Selector32~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector32~2_combout ),
	.cout());
defparam \Selector32~2 .lut_mask = 16'hFEFE;
defparam \Selector32~2 .sum_lutc_input = "datac";

dffeas \m_state.100000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector32~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.100000000~q ),
	.prn(vcc));
defparam \m_state.100000000 .is_wysiwyg = "true";
defparam \m_state.100000000 .power_up = "low";

cycloneive_lcell_comb \pending~10 (
	.dataa(\pending~4_combout ),
	.datab(\pending~9_combout ),
	.datac(gnd),
	.datad(\active_cs_n~q ),
	.cin(gnd),
	.combout(\pending~10_combout ),
	.cout());
defparam \pending~10 .lut_mask = 16'hEEFF;
defparam \pending~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_next~19 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\refresh_request~q ),
	.datad(\pending~10_combout ),
	.cin(gnd),
	.combout(\m_next~19_combout ),
	.cout());
defparam \m_next~19 .lut_mask = 16'hFEFF;
defparam \m_next~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector29~0 (
	.dataa(\m_state.100000000~q ),
	.datab(entries_1),
	.datac(entries_0),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector29~0_combout ),
	.cout());
defparam \Selector29~0 .lut_mask = 16'hFEFF;
defparam \Selector29~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector29~1 (
	.dataa(\m_state.000100000~q ),
	.datab(\LessThan1~0_combout ),
	.datac(\Selector29~0_combout ),
	.datad(\pending~10_combout ),
	.cin(gnd),
	.combout(\Selector29~1_combout ),
	.cout());
defparam \Selector29~1 .lut_mask = 16'hFEFF;
defparam \Selector29~1 .sum_lutc_input = "datac";

dffeas \m_state.000100000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector29~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000100000~q ),
	.prn(vcc));
defparam \m_state.000100000 .is_wysiwyg = "true";
defparam \m_state.000100000 .power_up = "low";

cycloneive_lcell_comb \Selector39~2 (
	.dataa(\m_state.000100000~q ),
	.datab(\m_state.000000100~q ),
	.datac(\LessThan1~0_combout ),
	.datad(\m_count[0]~q ),
	.cin(gnd),
	.combout(\Selector39~2_combout ),
	.cout());
defparam \Selector39~2 .lut_mask = 16'hEFFE;
defparam \Selector39~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~3 (
	.dataa(\m_count[0]~q ),
	.datab(\init_done~q ),
	.datac(\refresh_request~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector39~3_combout ),
	.cout());
defparam \Selector39~3 .lut_mask = 16'hFEFF;
defparam \Selector39~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~4 (
	.dataa(\m_state.010000000~q ),
	.datab(\Selector39~3_combout ),
	.datac(\m_state.001000000~q ),
	.datad(\m_count[0]~q ),
	.cin(gnd),
	.combout(\Selector39~4_combout ),
	.cout());
defparam \Selector39~4 .lut_mask = 16'hFFFE;
defparam \Selector39~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~5 (
	.dataa(\Selector39~2_combout ),
	.datab(\Selector39~4_combout ),
	.datac(\Selector39~7_combout ),
	.datad(\m_count[0]~q ),
	.cin(gnd),
	.combout(\Selector39~5_combout ),
	.cout());
defparam \Selector39~5 .lut_mask = 16'hFFFE;
defparam \Selector39~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~6 (
	.dataa(\Selector39~5_combout ),
	.datab(\m_state.100000000~q ),
	.datac(\m_next~19_combout ),
	.datad(\m_count[0]~q ),
	.cin(gnd),
	.combout(\Selector39~6_combout ),
	.cout());
defparam \Selector39~6 .lut_mask = 16'hFFFE;
defparam \Selector39~6 .sum_lutc_input = "datac";

dffeas \m_count[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector39~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_count[0]~q ),
	.prn(vcc));
defparam \m_count[0] .is_wysiwyg = "true";
defparam \m_count[0] .power_up = "low";

cycloneive_lcell_comb \m_count~0 (
	.dataa(\m_count[1]~q ),
	.datab(\m_count[0]~q ),
	.datac(\m_count[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\m_count~0_combout ),
	.cout());
defparam \m_count~0 .lut_mask = 16'hF6F6;
defparam \m_count~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~0 (
	.dataa(\m_count~0_combout ),
	.datab(gnd),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\Selector38~0_combout ),
	.cout());
defparam \Selector38~0 .lut_mask = 16'hAFFF;
defparam \Selector38~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~1 (
	.dataa(\m_state.000000001~q ),
	.datab(\m_count[1]~q ),
	.datac(\init_done~q ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector38~1_combout ),
	.cout());
defparam \Selector38~1 .lut_mask = 16'hEFFF;
defparam \Selector38~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~2 (
	.dataa(\Selector38~0_combout ),
	.datab(\Selector38~1_combout ),
	.datac(\m_count[1]~q ),
	.datad(\m_state.001000000~q ),
	.cin(gnd),
	.combout(\Selector38~2_combout ),
	.cout());
defparam \Selector38~2 .lut_mask = 16'hFEFF;
defparam \Selector38~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~3 (
	.dataa(\Selector38~2_combout ),
	.datab(\m_count[1]~q ),
	.datac(\m_next~19_combout ),
	.datad(\m_state.100000000~q ),
	.cin(gnd),
	.combout(\Selector38~3_combout ),
	.cout());
defparam \Selector38~3 .lut_mask = 16'hEFFF;
defparam \Selector38~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~4 (
	.dataa(gnd),
	.datab(\Selector41~0_combout ),
	.datac(\refresh_request~q ),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector38~4_combout ),
	.cout());
defparam \Selector38~4 .lut_mask = 16'h3FFF;
defparam \Selector38~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~5 (
	.dataa(\Selector38~3_combout ),
	.datab(\m_state.000001000~q ),
	.datac(\m_state.000010000~q ),
	.datad(\Selector38~4_combout ),
	.cin(gnd),
	.combout(\Selector38~5_combout ),
	.cout());
defparam \Selector38~5 .lut_mask = 16'hBFFF;
defparam \Selector38~5 .sum_lutc_input = "datac";

dffeas \m_count[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector38~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_count[1]~q ),
	.prn(vcc));
defparam \m_count[1] .is_wysiwyg = "true";
defparam \m_count[1] .power_up = "low";

cycloneive_lcell_comb \LessThan1~0 (
	.dataa(\m_count[2]~q ),
	.datab(\m_count[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan1~0_combout ),
	.cout());
defparam \LessThan1~0 .lut_mask = 16'hEEEE;
defparam \LessThan1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~0 (
	.dataa(\m_state.000000100~q ),
	.datab(\Selector32~0_combout ),
	.datac(\m_state.100000000~q ),
	.datad(\LessThan1~0_combout ),
	.cin(gnd),
	.combout(\Selector27~0_combout ),
	.cout());
defparam \Selector27~0 .lut_mask = 16'hEFFF;
defparam \Selector27~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector35~0 (
	.dataa(\active_rnw~q ),
	.datab(\m_state.010000000~q ),
	.datac(\m_state.100000000~q ),
	.datad(\m_next~19_combout ),
	.cin(gnd),
	.combout(\Selector35~0_combout ),
	.cout());
defparam \Selector35~0 .lut_mask = 16'h7FFF;
defparam \Selector35~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector25~4 (
	.dataa(\init_done~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector25~4_combout ),
	.cout());
defparam \Selector25~4 .lut_mask = 16'hAAFF;
defparam \Selector25~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector25~5 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\Selector25~4_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector25~5_combout ),
	.cout());
defparam \Selector25~5 .lut_mask = 16'hFEFF;
defparam \Selector25~5 .sum_lutc_input = "datac";

dffeas \m_state.000000010 (
	.clk(wire_pll7_clk_0),
	.d(\Selector25~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000010~q ),
	.prn(vcc));
defparam \m_state.000000010 .is_wysiwyg = "true";
defparam \m_state.000000010 .power_up = "low";

cycloneive_lcell_comb \Selector34~1 (
	.dataa(\m_state.000000010~q ),
	.datab(\m_state.010000000~q ),
	.datac(\m_state.100000000~q ),
	.datad(\m_next~19_combout ),
	.cin(gnd),
	.combout(\Selector34~1_combout ),
	.cout());
defparam \Selector34~1 .lut_mask = 16'hFFFE;
defparam \Selector34~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector34~2 (
	.dataa(\refresh_request~q ),
	.datab(\init_done~q ),
	.datac(\m_state.000000001~q ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector34~2_combout ),
	.cout());
defparam \Selector34~2 .lut_mask = 16'hDEFF;
defparam \Selector34~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector34~3 (
	.dataa(\Selector41~0_combout ),
	.datab(\Selector34~1_combout ),
	.datac(\m_state.000000001~q ),
	.datad(\Selector34~2_combout ),
	.cin(gnd),
	.combout(\Selector34~3_combout ),
	.cout());
defparam \Selector34~3 .lut_mask = 16'hEFFE;
defparam \Selector34~3 .sum_lutc_input = "datac";

dffeas \m_next.000010000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector35~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\m_state.000000010~q ),
	.sload(gnd),
	.ena(\Selector34~3_combout ),
	.q(\m_next.000010000~q ),
	.prn(vcc));
defparam \m_next.000010000 .is_wysiwyg = "true";
defparam \m_next.000010000 .power_up = "low";

cycloneive_lcell_comb \Selector27~1 (
	.dataa(\pending~10_combout ),
	.datab(\m_state.100000000~q ),
	.datac(\refresh_request~q ),
	.datad(\Selector32~0_combout ),
	.cin(gnd),
	.combout(\Selector27~1_combout ),
	.cout());
defparam \Selector27~1 .lut_mask = 16'hEFFF;
defparam \Selector27~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector28~0 (
	.dataa(\Selector27~0_combout ),
	.datab(\m_next.000010000~q ),
	.datac(\Selector27~1_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[42]~1_combout ),
	.cin(gnd),
	.combout(\Selector28~0_combout ),
	.cout());
defparam \Selector28~0 .lut_mask = 16'hFEFF;
defparam \Selector28~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~3 (
	.dataa(\refresh_request~q ),
	.datab(\m_state.000000001~q ),
	.datac(\Selector41~0_combout ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector27~3_combout ),
	.cout());
defparam \Selector27~3 .lut_mask = 16'hEFFF;
defparam \Selector27~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~4 (
	.dataa(\the_niosII_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(\refresh_request~q ),
	.datac(\init_done~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector27~4_combout ),
	.cout());
defparam \Selector27~4 .lut_mask = 16'hEFFF;
defparam \Selector27~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~5 (
	.dataa(\m_state.100000000~q ),
	.datab(\m_state.000000100~q ),
	.datac(\Selector32~0_combout ),
	.datad(\LessThan1~0_combout ),
	.cin(gnd),
	.combout(\Selector27~5_combout ),
	.cout());
defparam \Selector27~5 .lut_mask = 16'hEFFF;
defparam \Selector27~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr8~0 (
	.dataa(gnd),
	.datab(\m_state.000000010~q ),
	.datac(\m_state.001000000~q ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\WideOr8~0_combout ),
	.cout());
defparam \WideOr8~0 .lut_mask = 16'h3FFF;
defparam \WideOr8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~6 (
	.dataa(\Selector27~3_combout ),
	.datab(\Selector27~4_combout ),
	.datac(\Selector27~5_combout ),
	.datad(\WideOr8~0_combout ),
	.cin(gnd),
	.combout(\Selector27~6_combout ),
	.cout());
defparam \Selector27~6 .lut_mask = 16'hFEFF;
defparam \Selector27~6 .sum_lutc_input = "datac";

dffeas \m_state.000010000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector28~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector27~6_combout ),
	.q(\m_state.000010000~q ),
	.prn(vcc));
defparam \m_state.000010000 .is_wysiwyg = "true";
defparam \m_state.000010000 .power_up = "low";

cycloneive_lcell_comb \Selector39~7 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\Selector41~0_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector39~7_combout ),
	.cout());
defparam \Selector39~7 .lut_mask = 16'hEFFF;
defparam \Selector39~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector37~0 (
	.dataa(\m_state.000000100~q ),
	.datab(\m_state.000100000~q ),
	.datac(\m_count[1]~q ),
	.datad(\m_count[0]~q ),
	.cin(gnd),
	.combout(\Selector37~0_combout ),
	.cout());
defparam \Selector37~0 .lut_mask = 16'hFFFE;
defparam \Selector37~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector37~1 (
	.dataa(\init_done~q ),
	.datab(\refresh_request~q ),
	.datac(\m_state.000000001~q ),
	.datad(\m_state.001000000~q ),
	.cin(gnd),
	.combout(\Selector37~1_combout ),
	.cout());
defparam \Selector37~1 .lut_mask = 16'hFEFF;
defparam \Selector37~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector37~2 (
	.dataa(\Selector37~0_combout ),
	.datab(\m_next~19_combout ),
	.datac(\m_state.100000000~q ),
	.datad(\Selector37~1_combout ),
	.cin(gnd),
	.combout(\Selector37~2_combout ),
	.cout());
defparam \Selector37~2 .lut_mask = 16'hFFDF;
defparam \Selector37~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector37~3 (
	.dataa(\m_count[2]~q ),
	.datab(\m_state.010000000~q ),
	.datac(\Selector39~7_combout ),
	.datad(\Selector37~2_combout ),
	.cin(gnd),
	.combout(\Selector37~3_combout ),
	.cout());
defparam \Selector37~3 .lut_mask = 16'hFEFF;
defparam \Selector37~3 .sum_lutc_input = "datac";

dffeas \m_count[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector37~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_count[2]~q ),
	.prn(vcc));
defparam \m_count[2] .is_wysiwyg = "true";
defparam \m_count[2] .power_up = "low";

cycloneive_lcell_comb \Selector30~3 (
	.dataa(\m_count[2]~q ),
	.datab(\m_count[1]~q ),
	.datac(\Selector30~2_combout ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\Selector30~3_combout ),
	.cout());
defparam \Selector30~3 .lut_mask = 16'hFFF7;
defparam \Selector30~3 .sum_lutc_input = "datac";

dffeas \m_state.001000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector30~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.001000000~q ),
	.prn(vcc));
defparam \m_state.001000000 .is_wysiwyg = "true";
defparam \m_state.001000000 .power_up = "low";

cycloneive_lcell_comb \Selector36~0 (
	.dataa(\m_state.000000100~q ),
	.datab(\m_state.000100000~q ),
	.datac(\init_done~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector36~0_combout ),
	.cout());
defparam \Selector36~0 .lut_mask = 16'hFEFF;
defparam \Selector36~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector36~1 (
	.dataa(\m_state.001000000~q ),
	.datab(\Selector36~0_combout ),
	.datac(\m_state.100000000~q ),
	.datad(\m_next~19_combout ),
	.cin(gnd),
	.combout(\Selector36~1_combout ),
	.cout());
defparam \Selector36~1 .lut_mask = 16'hFEFF;
defparam \Selector36~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector36~2 (
	.dataa(\Selector30~2_combout ),
	.datab(\m_next.010000000~q ),
	.datac(\Selector36~1_combout ),
	.datad(\Selector39~7_combout ),
	.cin(gnd),
	.combout(\Selector36~2_combout ),
	.cout());
defparam \Selector36~2 .lut_mask = 16'hFFFE;
defparam \Selector36~2 .sum_lutc_input = "datac";

dffeas \m_next.010000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector36~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.010000000~q ),
	.prn(vcc));
defparam \m_next.010000000 .is_wysiwyg = "true";
defparam \m_next.010000000 .power_up = "low";

cycloneive_lcell_comb \Selector31~0 (
	.dataa(\m_state.000000100~q ),
	.datab(\m_next.010000000~q ),
	.datac(\m_count[2]~q ),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector31~0_combout ),
	.cout());
defparam \Selector31~0 .lut_mask = 16'hEFFF;
defparam \Selector31~0 .sum_lutc_input = "datac";

dffeas \m_state.010000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector31~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.010000000~q ),
	.prn(vcc));
defparam \m_state.010000000 .is_wysiwyg = "true";
defparam \m_state.010000000 .power_up = "low";

cycloneive_lcell_comb \Selector34~0 (
	.dataa(\active_rnw~q ),
	.datab(\m_state.100000000~q ),
	.datac(\m_next~19_combout ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\Selector34~0_combout ),
	.cout());
defparam \Selector34~0 .lut_mask = 16'hBFFF;
defparam \Selector34~0 .sum_lutc_input = "datac";

dffeas \m_next.000001000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector34~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\m_state.000000010~q ),
	.sload(gnd),
	.ena(\Selector34~3_combout ),
	.q(\m_next.000001000~q ),
	.prn(vcc));
defparam \m_next.000001000 .is_wysiwyg = "true";
defparam \m_next.000001000 .power_up = "low";

cycloneive_lcell_comb \Selector27~2 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[42]~1_combout ),
	.datab(\m_next.000001000~q ),
	.datac(\Selector27~0_combout ),
	.datad(\Selector27~1_combout ),
	.cin(gnd),
	.combout(\Selector27~2_combout ),
	.cout());
defparam \Selector27~2 .lut_mask = 16'hFFFE;
defparam \Selector27~2 .sum_lutc_input = "datac";

dffeas \m_state.000001000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector27~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector27~6_combout ),
	.q(\m_state.000001000~q ),
	.prn(vcc));
defparam \m_state.000001000 .is_wysiwyg = "true";
defparam \m_state.000001000 .power_up = "low";

cycloneive_lcell_comb \WideOr9~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\m_state.000001000~q ),
	.datad(\m_state.000010000~q ),
	.cin(gnd),
	.combout(\WideOr9~0_combout ),
	.cout());
defparam \WideOr9~0 .lut_mask = 16'h0FFF;
defparam \WideOr9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector26~0 (
	.dataa(\Selector41~0_combout ),
	.datab(\m_state.000000100~q ),
	.datac(\refresh_request~q ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
defparam \Selector26~0 .lut_mask = 16'hFEFF;
defparam \Selector26~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector26~1 (
	.dataa(\m_state.100000000~q ),
	.datab(\refresh_request~q ),
	.datac(gnd),
	.datad(\WideOr8~0_combout ),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
defparam \Selector26~1 .lut_mask = 16'hEEFF;
defparam \Selector26~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector26~2 (
	.dataa(\Selector26~0_combout ),
	.datab(\Selector26~1_combout ),
	.datac(\m_state.000000100~q ),
	.datad(\LessThan1~0_combout ),
	.cin(gnd),
	.combout(\Selector26~2_combout ),
	.cout());
defparam \Selector26~2 .lut_mask = 16'hFFFE;
defparam \Selector26~2 .sum_lutc_input = "datac";

dffeas \m_state.000000100 (
	.clk(wire_pll7_clk_0),
	.d(\Selector26~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000100~q ),
	.prn(vcc));
defparam \m_state.000000100 .is_wysiwyg = "true";
defparam \m_state.000000100 .power_up = "low";

cycloneive_lcell_comb \Selector33~0 (
	.dataa(\Selector41~0_combout ),
	.datab(\refresh_request~q ),
	.datac(\m_next.000000001~q ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector33~0_combout ),
	.cout());
defparam \Selector33~0 .lut_mask = 16'hEFFF;
defparam \Selector33~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_addr[1]~3 (
	.dataa(gnd),
	.datab(\m_state.100000000~q ),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\m_addr[1]~3_combout ),
	.cout());
defparam \m_addr[1]~3 .lut_mask = 16'h3FFF;
defparam \m_addr[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~1 (
	.dataa(\m_state.001000000~q ),
	.datab(\m_state.000000001~q ),
	.datac(\refresh_request~q ),
	.datad(\m_addr[1]~3_combout ),
	.cin(gnd),
	.combout(\Selector33~1_combout ),
	.cout());
defparam \Selector33~1 .lut_mask = 16'hBFFF;
defparam \Selector33~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~2 (
	.dataa(\Selector33~1_combout ),
	.datab(\init_done~q ),
	.datac(\m_state.000000001~q ),
	.datad(\m_next.000000001~q ),
	.cin(gnd),
	.combout(\Selector33~2_combout ),
	.cout());
defparam \Selector33~2 .lut_mask = 16'hFFFD;
defparam \Selector33~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~3 (
	.dataa(\m_state.100000000~q ),
	.datab(\refresh_request~q ),
	.datac(\the_niosII_sdram_input_efifo_module|Equal1~0_combout ),
	.datad(\pending~10_combout ),
	.cin(gnd),
	.combout(\Selector33~3_combout ),
	.cout());
defparam \Selector33~3 .lut_mask = 16'hFEFF;
defparam \Selector33~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~4 (
	.dataa(\m_state.010000000~q ),
	.datab(\Selector33~0_combout ),
	.datac(\Selector33~2_combout ),
	.datad(\Selector33~3_combout ),
	.cin(gnd),
	.combout(\Selector33~4_combout ),
	.cout());
defparam \Selector33~4 .lut_mask = 16'hF7FF;
defparam \Selector33~4 .sum_lutc_input = "datac";

dffeas \m_next.000000001 (
	.clk(wire_pll7_clk_0),
	.d(\Selector33~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.000000001~q ),
	.prn(vcc));
defparam \m_next.000000001 .is_wysiwyg = "true";
defparam \m_next.000000001 .power_up = "low";

cycloneive_lcell_comb \Selector24~0 (
	.dataa(\m_state.000000100~q ),
	.datab(\m_count[2]~q ),
	.datac(\m_count[1]~q ),
	.datad(\m_next.000000001~q ),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
defparam \Selector24~0 .lut_mask = 16'hBFFF;
defparam \Selector24~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector24~1 (
	.dataa(\Selector24~0_combout ),
	.datab(\Selector32~0_combout ),
	.datac(\init_done~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector24~1_combout ),
	.cout());
defparam \Selector24~1 .lut_mask = 16'hFFF7;
defparam \Selector24~1 .sum_lutc_input = "datac";

dffeas \m_state.000000001 (
	.clk(wire_pll7_clk_0),
	.d(\Selector24~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000001~q ),
	.prn(vcc));
defparam \m_state.000000001 .is_wysiwyg = "true";
defparam \m_state.000000001 .power_up = "low";

cycloneive_lcell_comb \Selector23~0 (
	.dataa(\m_state.000000001~q ),
	.datab(\ack_refresh_request~q ),
	.datac(\m_state.010000000~q ),
	.datad(\init_done~q ),
	.cin(gnd),
	.combout(\Selector23~0_combout ),
	.cout());
defparam \Selector23~0 .lut_mask = 16'hFEFF;
defparam \Selector23~0 .sum_lutc_input = "datac";

dffeas ack_refresh_request(
	.clk(wire_pll7_clk_0),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ack_refresh_request~q ),
	.prn(vcc));
defparam ack_refresh_request.is_wysiwyg = "true";
defparam ack_refresh_request.power_up = "low";

cycloneive_lcell_comb \refresh_request~0 (
	.dataa(\init_done~q ),
	.datab(\refresh_request~q ),
	.datac(\Equal0~4_combout ),
	.datad(\ack_refresh_request~q ),
	.cin(gnd),
	.combout(\refresh_request~0_combout ),
	.cout());
defparam \refresh_request~0 .lut_mask = 16'hFEFF;
defparam \refresh_request~0 .sum_lutc_input = "datac";

dffeas refresh_request(
	.clk(wire_pll7_clk_0),
	.d(\refresh_request~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_request~q ),
	.prn(vcc));
defparam refresh_request.is_wysiwyg = "true";
defparam refresh_request.power_up = "low";

cycloneive_lcell_comb \active_rnw~0 (
	.dataa(\m_state.000000001~q ),
	.datab(\the_niosII_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(\init_done~q ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\active_rnw~0_combout ),
	.cout());
defparam \active_rnw~0 .lut_mask = 16'hFFD8;
defparam \active_rnw~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_rnw~1 (
	.dataa(\m_state.100000000~q ),
	.datab(\Selector41~0_combout ),
	.datac(\m_state.000000001~q ),
	.datad(\active_rnw~0_combout ),
	.cin(gnd),
	.combout(\active_rnw~1_combout ),
	.cout());
defparam \active_rnw~1 .lut_mask = 16'hEFFE;
defparam \active_rnw~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_rnw~2 (
	.dataa(r_sync_rst),
	.datab(\refresh_request~q ),
	.datac(\active_rnw~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\active_rnw~2_combout ),
	.cout());
defparam \active_rnw~2 .lut_mask = 16'hF7F7;
defparam \active_rnw~2 .sum_lutc_input = "datac";

dffeas \active_addr[10] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[28]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[10]~q ),
	.prn(vcc));
defparam \active_addr[10] .is_wysiwyg = "true";
defparam \active_addr[10] .power_up = "low";

cycloneive_lcell_comb \Selector41~1 (
	.dataa(\Selector41~0_combout ),
	.datab(\m_state.100000000~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector41~1_combout ),
	.cout());
defparam \Selector41~1 .lut_mask = 16'hEFFF;
defparam \Selector41~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector41~2 (
	.dataa(\Selector41~1_combout ),
	.datab(\the_niosII_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(\Selector25~4_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector41~2_combout ),
	.cout());
defparam \Selector41~2 .lut_mask = 16'hFEFF;
defparam \Selector41~2 .sum_lutc_input = "datac";

dffeas f_pop(
	.clk(wire_pll7_clk_0),
	.d(\Selector41~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\f_pop~q ),
	.prn(vcc));
defparam f_pop.is_wysiwyg = "true";
defparam f_pop.power_up = "low";

cycloneive_lcell_comb \m_addr[1]~2 (
	.dataa(\m_state.000000010~q ),
	.datab(\f_pop~q ),
	.datac(\Selector41~0_combout ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\m_addr[1]~2_combout ),
	.cout());
defparam \m_addr[1]~2 .lut_mask = 16'hFAFC;
defparam \m_addr[1]~2 .sum_lutc_input = "datac";

dffeas \active_addr[0] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[18]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[0]~q ),
	.prn(vcc));
defparam \active_addr[0] .is_wysiwyg = "true";
defparam \active_addr[0] .power_up = "low";

dffeas \i_addr[12] (
	.clk(wire_pll7_clk_0),
	.d(\i_state.111~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_addr[12]~q ),
	.prn(vcc));
defparam \i_addr[12] .is_wysiwyg = "true";
defparam \i_addr[12] .power_up = "low";

cycloneive_lcell_comb \Selector97~0 (
	.dataa(\m_addr[1]~2_combout ),
	.datab(\active_addr[0]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector97~0_combout ),
	.cout());
defparam \Selector97~0 .lut_mask = 16'hDEFF;
defparam \Selector97~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector97~1 (
	.dataa(\active_addr[10]~q ),
	.datab(\m_addr[1]~2_combout ),
	.datac(\Selector97~0_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[18]~16_combout ),
	.cin(gnd),
	.combout(\Selector97~1_combout ),
	.cout());
defparam \Selector97~1 .lut_mask = 16'hFFBE;
defparam \Selector97~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_addr[1]~4 (
	.dataa(\init_done~q ),
	.datab(\m_state.000000001~q ),
	.datac(\m_state.010000000~q ),
	.datad(\m_addr[1]~3_combout ),
	.cin(gnd),
	.combout(\m_addr[1]~4_combout ),
	.cout());
defparam \m_addr[1]~4 .lut_mask = 16'hFFDF;
defparam \m_addr[1]~4 .sum_lutc_input = "datac";

dffeas \active_addr[1] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[19]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[1]~q ),
	.prn(vcc));
defparam \active_addr[1] .is_wysiwyg = "true";
defparam \active_addr[1] .power_up = "low";

cycloneive_lcell_comb \Selector96~0 (
	.dataa(\m_addr[1]~2_combout ),
	.datab(\active_addr[1]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector96~0_combout ),
	.cout());
defparam \Selector96~0 .lut_mask = 16'hDEFF;
defparam \Selector96~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector96~1 (
	.dataa(\active_addr[11]~q ),
	.datab(\m_addr[1]~2_combout ),
	.datac(\Selector96~0_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[19]~17_combout ),
	.cin(gnd),
	.combout(\Selector96~1_combout ),
	.cout());
defparam \Selector96~1 .lut_mask = 16'hFFBE;
defparam \Selector96~1 .sum_lutc_input = "datac";

dffeas \active_addr[2] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[20]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[2]~q ),
	.prn(vcc));
defparam \active_addr[2] .is_wysiwyg = "true";
defparam \active_addr[2] .power_up = "low";

cycloneive_lcell_comb \Selector95~0 (
	.dataa(\m_addr[1]~2_combout ),
	.datab(\active_addr[2]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector95~0_combout ),
	.cout());
defparam \Selector95~0 .lut_mask = 16'hDEFF;
defparam \Selector95~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector95~1 (
	.dataa(\active_addr[12]~q ),
	.datab(\m_addr[1]~2_combout ),
	.datac(\Selector95~0_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[20]~18_combout ),
	.cin(gnd),
	.combout(\Selector95~1_combout ),
	.cout());
defparam \Selector95~1 .lut_mask = 16'hFFBE;
defparam \Selector95~1 .sum_lutc_input = "datac";

dffeas \active_addr[3] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[21]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[3]~q ),
	.prn(vcc));
defparam \active_addr[3] .is_wysiwyg = "true";
defparam \active_addr[3] .power_up = "low";

cycloneive_lcell_comb \Selector94~0 (
	.dataa(\m_addr[1]~2_combout ),
	.datab(\active_addr[3]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector94~0_combout ),
	.cout());
defparam \Selector94~0 .lut_mask = 16'hDEFF;
defparam \Selector94~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector94~1 (
	.dataa(\active_addr[13]~q ),
	.datab(\m_addr[1]~2_combout ),
	.datac(\Selector94~0_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[21]~19_combout ),
	.cin(gnd),
	.combout(\Selector94~1_combout ),
	.cout());
defparam \Selector94~1 .lut_mask = 16'hFFBE;
defparam \Selector94~1 .sum_lutc_input = "datac";

dffeas \active_addr[4] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[22]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[4]~q ),
	.prn(vcc));
defparam \active_addr[4] .is_wysiwyg = "true";
defparam \active_addr[4] .power_up = "low";

cycloneive_lcell_comb \Selector93~0 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[22]~20_combout ),
	.datab(\active_addr[4]~q ),
	.datac(\f_pop~q ),
	.datad(\Selector41~0_combout ),
	.cin(gnd),
	.combout(\Selector93~0_combout ),
	.cout());
defparam \Selector93~0 .lut_mask = 16'hEFFE;
defparam \Selector93~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector93~1 (
	.dataa(\active_addr[14]~q ),
	.datab(\Selector93~0_combout ),
	.datac(\WideOr9~0_combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector93~1_combout ),
	.cout());
defparam \Selector93~1 .lut_mask = 16'hACFF;
defparam \Selector93~1 .sum_lutc_input = "datac";

dffeas \active_addr[5] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[23]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[5]~q ),
	.prn(vcc));
defparam \active_addr[5] .is_wysiwyg = "true";
defparam \active_addr[5] .power_up = "low";

cycloneive_lcell_comb f_select(
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\f_pop~q ),
	.datad(\pending~10_combout ),
	.cin(gnd),
	.combout(\f_select~combout ),
	.cout());
defparam f_select.lut_mask = 16'hFFFE;
defparam f_select.sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector92~0 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[23]~21_combout ),
	.datab(\active_addr[5]~q ),
	.datac(\f_select~combout ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector92~0_combout ),
	.cout());
defparam \Selector92~0 .lut_mask = 16'hACFF;
defparam \Selector92~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector92~1 (
	.dataa(\Selector92~0_combout ),
	.datab(\WideOr9~0_combout ),
	.datac(\active_addr[15]~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector92~1_combout ),
	.cout());
defparam \Selector92~1 .lut_mask = 16'hFEFF;
defparam \Selector92~1 .sum_lutc_input = "datac";

dffeas \active_addr[6] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[24]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[6]~q ),
	.prn(vcc));
defparam \active_addr[6] .is_wysiwyg = "true";
defparam \active_addr[6] .power_up = "low";

cycloneive_lcell_comb \Selector91~0 (
	.dataa(\m_addr[1]~2_combout ),
	.datab(\active_addr[6]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector91~0_combout ),
	.cout());
defparam \Selector91~0 .lut_mask = 16'hDEFF;
defparam \Selector91~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector91~1 (
	.dataa(\active_addr[16]~q ),
	.datab(\m_addr[1]~2_combout ),
	.datac(\Selector91~0_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[24]~22_combout ),
	.cin(gnd),
	.combout(\Selector91~1_combout ),
	.cout());
defparam \Selector91~1 .lut_mask = 16'hFFBE;
defparam \Selector91~1 .sum_lutc_input = "datac";

dffeas \active_addr[7] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[25]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[7]~q ),
	.prn(vcc));
defparam \active_addr[7] .is_wysiwyg = "true";
defparam \active_addr[7] .power_up = "low";

cycloneive_lcell_comb \Selector90~0 (
	.dataa(\m_addr[1]~2_combout ),
	.datab(\active_addr[7]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector90~0_combout ),
	.cout());
defparam \Selector90~0 .lut_mask = 16'hDEFF;
defparam \Selector90~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector90~1 (
	.dataa(\active_addr[17]~q ),
	.datab(\m_addr[1]~2_combout ),
	.datac(\Selector90~0_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[25]~23_combout ),
	.cin(gnd),
	.combout(\Selector90~1_combout ),
	.cout());
defparam \Selector90~1 .lut_mask = 16'hFFBE;
defparam \Selector90~1 .sum_lutc_input = "datac";

dffeas \active_addr[8] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[26]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_addr[8]~q ),
	.prn(vcc));
defparam \active_addr[8] .is_wysiwyg = "true";
defparam \active_addr[8] .power_up = "low";

cycloneive_lcell_comb \Selector89~0 (
	.dataa(\m_addr[1]~2_combout ),
	.datab(\active_addr[8]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector89~0_combout ),
	.cout());
defparam \Selector89~0 .lut_mask = 16'hDEFF;
defparam \Selector89~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector89~1 (
	.dataa(\active_addr[18]~q ),
	.datab(\m_addr[1]~2_combout ),
	.datac(\Selector89~0_combout ),
	.datad(\the_niosII_sdram_input_efifo_module|rd_data[26]~24_combout ),
	.cin(gnd),
	.combout(\Selector89~1_combout ),
	.cout());
defparam \Selector89~1 .lut_mask = 16'hFFBE;
defparam \Selector89~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always5~0 (
	.dataa(\f_pop~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Selector41~0_combout ),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'hFF55;
defparam \always5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector88~2 (
	.dataa(\active_addr[19]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector88~2_combout ),
	.cout());
defparam \Selector88~2 .lut_mask = 16'h88BB;
defparam \Selector88~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector88~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector88~2_combout ),
	.cin(gnd),
	.combout(\Selector88~3_combout ),
	.cout());
defparam \Selector88~3 .lut_mask = 16'hFFF7;
defparam \Selector88~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector87~2 (
	.dataa(\active_addr[20]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector87~2_combout ),
	.cout());
defparam \Selector87~2 .lut_mask = 16'h88BB;
defparam \Selector87~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector87~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector87~2_combout ),
	.cin(gnd),
	.combout(\Selector87~3_combout ),
	.cout());
defparam \Selector87~3 .lut_mask = 16'hFFF7;
defparam \Selector87~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector86~2 (
	.dataa(\active_addr[21]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector86~2_combout ),
	.cout());
defparam \Selector86~2 .lut_mask = 16'h88BB;
defparam \Selector86~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector86~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector86~2_combout ),
	.cin(gnd),
	.combout(\Selector86~3_combout ),
	.cout());
defparam \Selector86~3 .lut_mask = 16'hFFF7;
defparam \Selector86~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector85~2 (
	.dataa(\active_addr[22]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector85~2_combout ),
	.cout());
defparam \Selector85~2 .lut_mask = 16'h88BB;
defparam \Selector85~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector85~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector85~2_combout ),
	.cin(gnd),
	.combout(\Selector85~3_combout ),
	.cout());
defparam \Selector85~3 .lut_mask = 16'hFFF7;
defparam \Selector85~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector99~0 (
	.dataa(\active_addr[9]~q ),
	.datab(\the_niosII_sdram_input_efifo_module|rd_data[27]~0_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector99~0_combout ),
	.cout());
defparam \Selector99~0 .lut_mask = 16'hEFFE;
defparam \Selector99~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr16~0 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.000000010~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr16~0_combout ),
	.cout());
defparam \WideOr16~0 .lut_mask = 16'hFEFE;
defparam \WideOr16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector98~0 (
	.dataa(\active_addr[23]~q ),
	.datab(\the_niosII_sdram_input_efifo_module|rd_data[41]~2_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector98~0_combout ),
	.cout());
defparam \Selector98~0 .lut_mask = 16'hEFFE;
defparam \Selector98~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\i_state.001~q ),
	.datab(\i_state.101~q ),
	.datac(\i_cmd[1]~q ),
	.datad(\WideOr6~0_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFFF7;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \i_cmd[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[1]~q ),
	.prn(vcc));
defparam \i_cmd[1] .is_wysiwyg = "true";
defparam \i_cmd[1] .power_up = "low";

cycloneive_lcell_comb \Selector21~0 (
	.dataa(\init_done~q ),
	.datab(\i_cmd[1]~q ),
	.datac(\m_state.000000001~q ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
defparam \Selector21~0 .lut_mask = 16'hDFD5;
defparam \Selector21~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector21~1 (
	.dataa(\always5~0_combout ),
	.datab(\WideOr9~0_combout ),
	.datac(\m_state.000000001~q ),
	.datad(\Selector21~0_combout ),
	.cin(gnd),
	.combout(\Selector21~1_combout ),
	.cout());
defparam \Selector21~1 .lut_mask = 16'hFFB8;
defparam \Selector21~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\i_state.101~q ),
	.datab(gnd),
	.datac(\i_cmd[3]~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hFFF5;
defparam \Selector0~0 .sum_lutc_input = "datac";

dffeas \i_cmd[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[3]~q ),
	.prn(vcc));
defparam \i_cmd[3] .is_wysiwyg = "true";
defparam \i_cmd[3] .power_up = "low";

cycloneive_lcell_comb \Selector19~0 (
	.dataa(\init_done~q ),
	.datab(\i_cmd[3]~q ),
	.datac(\refresh_request~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
defparam \Selector19~0 .lut_mask = 16'h27FF;
defparam \Selector19~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~1 (
	.dataa(\m_state.000000001~q ),
	.datab(\m_state.001000000~q ),
	.datac(\m_state.010000000~q ),
	.datad(\m_state.000000100~q ),
	.cin(gnd),
	.combout(\Selector19~1_combout ),
	.cout());
defparam \Selector19~1 .lut_mask = 16'hBFFF;
defparam \Selector19~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~2 (
	.dataa(\m_state.001000000~q ),
	.datab(\m_state.000000100~q ),
	.datac(\refresh_request~q ),
	.datad(\m_next.010000000~q ),
	.cin(gnd),
	.combout(\Selector19~2_combout ),
	.cout());
defparam \Selector19~2 .lut_mask = 16'hEFFF;
defparam \Selector19~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~3 (
	.dataa(\Selector19~0_combout ),
	.datab(\active_cs_n~q ),
	.datac(\Selector19~1_combout ),
	.datad(\Selector19~2_combout ),
	.cin(gnd),
	.combout(\Selector19~3_combout ),
	.cout());
defparam \Selector19~3 .lut_mask = 16'h7FFF;
defparam \Selector19~3 .sum_lutc_input = "datac";

dffeas \active_dqm[0] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[16]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_dqm[0]~q ),
	.prn(vcc));
defparam \active_dqm[0] .is_wysiwyg = "true";
defparam \active_dqm[0] .power_up = "low";

cycloneive_lcell_comb \Selector117~0 (
	.dataa(\active_dqm[0]~q ),
	.datab(\the_niosII_sdram_input_efifo_module|rd_data[16]~25_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector117~0_combout ),
	.cout());
defparam \Selector117~0 .lut_mask = 16'hEFFE;
defparam \Selector117~0 .sum_lutc_input = "datac";

dffeas \active_dqm[1] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[17]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_dqm[1]~q ),
	.prn(vcc));
defparam \active_dqm[1] .is_wysiwyg = "true";
defparam \active_dqm[1] .power_up = "low";

cycloneive_lcell_comb \Selector116~0 (
	.dataa(\active_dqm[1]~q ),
	.datab(\the_niosII_sdram_input_efifo_module|rd_data[17]~26_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector116~0_combout ),
	.cout());
defparam \Selector116~0 .lut_mask = 16'hEFFE;
defparam \Selector116~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_state.101~q ),
	.datac(\i_cmd[2]~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hFFF7;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \i_cmd[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[2]~q ),
	.prn(vcc));
defparam \i_cmd[2] .is_wysiwyg = "true";
defparam \i_cmd[2] .power_up = "low";

cycloneive_lcell_comb \Selector20~0 (
	.dataa(\WideOr8~0_combout ),
	.datab(\init_done~q ),
	.datac(\i_cmd[2]~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
defparam \Selector20~0 .lut_mask = 16'hF377;
defparam \Selector20~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\i_state.010~q ),
	.datab(\i_state.101~q ),
	.datac(\i_cmd[0]~q ),
	.datad(\WideOr6~0_combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hFFF7;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas \i_cmd[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[0]~q ),
	.prn(vcc));
defparam \i_cmd[0] .is_wysiwyg = "true";
defparam \i_cmd[0] .power_up = "low";

cycloneive_lcell_comb \Selector22~0 (
	.dataa(\init_done~q ),
	.datab(\i_cmd[0]~q ),
	.datac(\m_state.000000001~q ),
	.datad(\m_state.001000000~q ),
	.cin(gnd),
	.combout(\Selector22~0_combout ),
	.cout());
defparam \Selector22~0 .lut_mask = 16'hDFD5;
defparam \Selector22~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector22~1 (
	.dataa(\m_state.000010000~q ),
	.datab(\always5~0_combout ),
	.datac(\m_state.000000001~q ),
	.datad(\Selector22~0_combout ),
	.cin(gnd),
	.combout(\Selector22~1_combout ),
	.cout());
defparam \Selector22~1 .lut_mask = 16'hFFD8;
defparam \Selector22~1 .sum_lutc_input = "datac";

dffeas \active_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[0]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[0]~q ),
	.prn(vcc));
defparam \active_data[0] .is_wysiwyg = "true";
defparam \active_data[0] .power_up = "low";

cycloneive_lcell_comb \Selector115~0 (
	.dataa(\active_data[0]~q ),
	.datab(m_data_0),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector115~0_combout ),
	.cout());
defparam \Selector115~0 .lut_mask = 16'hEFFE;
defparam \Selector115~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_data[1]~0 (
	.dataa(\f_pop~q ),
	.datab(\Selector41~0_combout ),
	.datac(\m_state.000010000~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\m_data[1]~0_combout ),
	.cout());
defparam \m_data[1]~0 .lut_mask = 16'hFEFE;
defparam \m_data[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector115~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[0]~27_combout ),
	.datab(\Selector115~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector115~1_combout ),
	.cout());
defparam \Selector115~1 .lut_mask = 16'hAACC;
defparam \Selector115~1 .sum_lutc_input = "datac";

dffeas \active_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[1]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[1]~q ),
	.prn(vcc));
defparam \active_data[1] .is_wysiwyg = "true";
defparam \active_data[1] .power_up = "low";

cycloneive_lcell_comb \Selector114~0 (
	.dataa(\active_data[1]~q ),
	.datab(m_data_1),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector114~0_combout ),
	.cout());
defparam \Selector114~0 .lut_mask = 16'hEFFE;
defparam \Selector114~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector114~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[1]~28_combout ),
	.datab(\Selector114~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector114~1_combout ),
	.cout());
defparam \Selector114~1 .lut_mask = 16'hAACC;
defparam \Selector114~1 .sum_lutc_input = "datac";

dffeas \active_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[2]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[2]~q ),
	.prn(vcc));
defparam \active_data[2] .is_wysiwyg = "true";
defparam \active_data[2] .power_up = "low";

cycloneive_lcell_comb \Selector113~0 (
	.dataa(\active_data[2]~q ),
	.datab(m_data_2),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector113~0_combout ),
	.cout());
defparam \Selector113~0 .lut_mask = 16'hEFFE;
defparam \Selector113~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector113~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[2]~29_combout ),
	.datab(\Selector113~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector113~1_combout ),
	.cout());
defparam \Selector113~1 .lut_mask = 16'hAACC;
defparam \Selector113~1 .sum_lutc_input = "datac";

dffeas \active_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[3]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[3]~q ),
	.prn(vcc));
defparam \active_data[3] .is_wysiwyg = "true";
defparam \active_data[3] .power_up = "low";

cycloneive_lcell_comb \Selector112~0 (
	.dataa(\active_data[3]~q ),
	.datab(m_data_3),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector112~0_combout ),
	.cout());
defparam \Selector112~0 .lut_mask = 16'hEFFE;
defparam \Selector112~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector112~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[3]~30_combout ),
	.datab(\Selector112~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector112~1_combout ),
	.cout());
defparam \Selector112~1 .lut_mask = 16'hAACC;
defparam \Selector112~1 .sum_lutc_input = "datac";

dffeas \active_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[4]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[4]~q ),
	.prn(vcc));
defparam \active_data[4] .is_wysiwyg = "true";
defparam \active_data[4] .power_up = "low";

cycloneive_lcell_comb \Selector111~0 (
	.dataa(\active_data[4]~q ),
	.datab(m_data_4),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector111~0_combout ),
	.cout());
defparam \Selector111~0 .lut_mask = 16'hEFFE;
defparam \Selector111~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector111~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[4]~31_combout ),
	.datab(\Selector111~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector111~1_combout ),
	.cout());
defparam \Selector111~1 .lut_mask = 16'hAACC;
defparam \Selector111~1 .sum_lutc_input = "datac";

dffeas \active_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[5]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[5]~q ),
	.prn(vcc));
defparam \active_data[5] .is_wysiwyg = "true";
defparam \active_data[5] .power_up = "low";

cycloneive_lcell_comb \Selector110~0 (
	.dataa(\active_data[5]~q ),
	.datab(m_data_5),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector110~0_combout ),
	.cout());
defparam \Selector110~0 .lut_mask = 16'hEFFE;
defparam \Selector110~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector110~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[5]~32_combout ),
	.datab(\Selector110~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector110~1_combout ),
	.cout());
defparam \Selector110~1 .lut_mask = 16'hAACC;
defparam \Selector110~1 .sum_lutc_input = "datac";

dffeas \active_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[6]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[6]~q ),
	.prn(vcc));
defparam \active_data[6] .is_wysiwyg = "true";
defparam \active_data[6] .power_up = "low";

cycloneive_lcell_comb \Selector109~0 (
	.dataa(\active_data[6]~q ),
	.datab(m_data_6),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector109~0_combout ),
	.cout());
defparam \Selector109~0 .lut_mask = 16'hEFFE;
defparam \Selector109~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector109~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[6]~33_combout ),
	.datab(\Selector109~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector109~1_combout ),
	.cout());
defparam \Selector109~1 .lut_mask = 16'hAACC;
defparam \Selector109~1 .sum_lutc_input = "datac";

dffeas \active_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[7]~q ),
	.prn(vcc));
defparam \active_data[7] .is_wysiwyg = "true";
defparam \active_data[7] .power_up = "low";

cycloneive_lcell_comb \Selector108~0 (
	.dataa(\active_data[7]~q ),
	.datab(m_data_7),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector108~0_combout ),
	.cout());
defparam \Selector108~0 .lut_mask = 16'hEFFE;
defparam \Selector108~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector108~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[7]~34_combout ),
	.datab(\Selector108~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector108~1_combout ),
	.cout());
defparam \Selector108~1 .lut_mask = 16'hAACC;
defparam \Selector108~1 .sum_lutc_input = "datac";

dffeas \active_data[8] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[8]~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[8]~q ),
	.prn(vcc));
defparam \active_data[8] .is_wysiwyg = "true";
defparam \active_data[8] .power_up = "low";

cycloneive_lcell_comb \Selector107~0 (
	.dataa(\active_data[8]~q ),
	.datab(m_data_8),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector107~0_combout ),
	.cout());
defparam \Selector107~0 .lut_mask = 16'hEFFE;
defparam \Selector107~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector107~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[8]~35_combout ),
	.datab(\Selector107~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector107~1_combout ),
	.cout());
defparam \Selector107~1 .lut_mask = 16'hAACC;
defparam \Selector107~1 .sum_lutc_input = "datac";

dffeas \active_data[9] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[9]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[9]~q ),
	.prn(vcc));
defparam \active_data[9] .is_wysiwyg = "true";
defparam \active_data[9] .power_up = "low";

cycloneive_lcell_comb \Selector106~0 (
	.dataa(\active_data[9]~q ),
	.datab(m_data_9),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector106~0_combout ),
	.cout());
defparam \Selector106~0 .lut_mask = 16'hEFFE;
defparam \Selector106~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector106~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[9]~36_combout ),
	.datab(\Selector106~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector106~1_combout ),
	.cout());
defparam \Selector106~1 .lut_mask = 16'hAACC;
defparam \Selector106~1 .sum_lutc_input = "datac";

dffeas \active_data[10] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[10]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[10]~q ),
	.prn(vcc));
defparam \active_data[10] .is_wysiwyg = "true";
defparam \active_data[10] .power_up = "low";

cycloneive_lcell_comb \Selector105~0 (
	.dataa(\active_data[10]~q ),
	.datab(m_data_10),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector105~0_combout ),
	.cout());
defparam \Selector105~0 .lut_mask = 16'hEFFE;
defparam \Selector105~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector105~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[10]~37_combout ),
	.datab(\Selector105~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector105~1_combout ),
	.cout());
defparam \Selector105~1 .lut_mask = 16'hAACC;
defparam \Selector105~1 .sum_lutc_input = "datac";

dffeas \active_data[11] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[11]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[11]~q ),
	.prn(vcc));
defparam \active_data[11] .is_wysiwyg = "true";
defparam \active_data[11] .power_up = "low";

cycloneive_lcell_comb \Selector104~0 (
	.dataa(\active_data[11]~q ),
	.datab(m_data_11),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector104~0_combout ),
	.cout());
defparam \Selector104~0 .lut_mask = 16'hEFFE;
defparam \Selector104~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector104~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[11]~38_combout ),
	.datab(\Selector104~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector104~1_combout ),
	.cout());
defparam \Selector104~1 .lut_mask = 16'hAACC;
defparam \Selector104~1 .sum_lutc_input = "datac";

dffeas \active_data[12] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[12]~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[12]~q ),
	.prn(vcc));
defparam \active_data[12] .is_wysiwyg = "true";
defparam \active_data[12] .power_up = "low";

cycloneive_lcell_comb \Selector103~0 (
	.dataa(\active_data[12]~q ),
	.datab(m_data_12),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector103~0_combout ),
	.cout());
defparam \Selector103~0 .lut_mask = 16'hEFFE;
defparam \Selector103~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector103~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[12]~39_combout ),
	.datab(\Selector103~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector103~1_combout ),
	.cout());
defparam \Selector103~1 .lut_mask = 16'hAACC;
defparam \Selector103~1 .sum_lutc_input = "datac";

dffeas \active_data[13] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[13]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[13]~q ),
	.prn(vcc));
defparam \active_data[13] .is_wysiwyg = "true";
defparam \active_data[13] .power_up = "low";

cycloneive_lcell_comb \Selector102~0 (
	.dataa(\active_data[13]~q ),
	.datab(m_data_13),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector102~0_combout ),
	.cout());
defparam \Selector102~0 .lut_mask = 16'hEFFE;
defparam \Selector102~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector102~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[13]~40_combout ),
	.datab(\Selector102~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector102~1_combout ),
	.cout());
defparam \Selector102~1 .lut_mask = 16'hAACC;
defparam \Selector102~1 .sum_lutc_input = "datac";

dffeas \active_data[14] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[14]~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[14]~q ),
	.prn(vcc));
defparam \active_data[14] .is_wysiwyg = "true";
defparam \active_data[14] .power_up = "low";

cycloneive_lcell_comb \Selector101~0 (
	.dataa(\active_data[14]~q ),
	.datab(m_data_14),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector101~0_combout ),
	.cout());
defparam \Selector101~0 .lut_mask = 16'hEFFE;
defparam \Selector101~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector101~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[14]~41_combout ),
	.datab(\Selector101~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector101~1_combout ),
	.cout());
defparam \Selector101~1 .lut_mask = 16'hAACC;
defparam \Selector101~1 .sum_lutc_input = "datac";

dffeas \active_data[15] (
	.clk(wire_pll7_clk_0),
	.d(\the_niosII_sdram_input_efifo_module|rd_data[15]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~2_combout ),
	.q(\active_data[15]~q ),
	.prn(vcc));
defparam \active_data[15] .is_wysiwyg = "true";
defparam \active_data[15] .power_up = "low";

cycloneive_lcell_comb \Selector100~0 (
	.dataa(\active_data[15]~q ),
	.datab(m_data_15),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector100~0_combout ),
	.cout());
defparam \Selector100~0 .lut_mask = 16'hEFFE;
defparam \Selector100~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector100~1 (
	.dataa(\the_niosII_sdram_input_efifo_module|rd_data[15]~42_combout ),
	.datab(\Selector100~0_combout ),
	.datac(gnd),
	.datad(\m_data[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector100~1_combout ),
	.cout());
defparam \Selector100~1 .lut_mask = 16'hAACC;
defparam \Selector100~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal4~0 (
	.dataa(m_cmd_1),
	.datab(gnd),
	.datac(m_cmd_2),
	.datad(m_cmd_0),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'hAFFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

dffeas \rd_valid[0] (
	.clk(wire_pll7_clk_0),
	.d(\Equal4~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[0]~q ),
	.prn(vcc));
defparam \rd_valid[0] .is_wysiwyg = "true";
defparam \rd_valid[0] .power_up = "low";

dffeas \rd_valid[1] (
	.clk(wire_pll7_clk_0),
	.d(\rd_valid[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[1]~q ),
	.prn(vcc));
defparam \rd_valid[1] .is_wysiwyg = "true";
defparam \rd_valid[1] .power_up = "low";

dffeas \rd_valid[2] (
	.clk(wire_pll7_clk_0),
	.d(\rd_valid[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[2]~q ),
	.prn(vcc));
defparam \rd_valid[2] .is_wysiwyg = "true";
defparam \rd_valid[2] .power_up = "low";

endmodule

module niosII_niosII_sdram_input_efifo_module (
	clk,
	reset_n,
	f_pop,
	entries_1,
	entries_0,
	Equal1,
	rd_data_27,
	rd_data_42,
	rd_data_41,
	rd_data_28,
	rd_data_30,
	rd_data_29,
	rd_data_32,
	rd_data_31,
	rd_data_34,
	rd_data_33,
	rd_data_36,
	rd_data_35,
	rd_data_38,
	rd_data_37,
	rd_data_40,
	rd_data_39,
	Selector41,
	rd_data_18,
	rd_data_19,
	rd_data_20,
	rd_data_21,
	rd_data_22,
	rd_data_23,
	rd_data_24,
	rd_data_25,
	rd_data_26,
	rd_data_16,
	rd_data_17,
	saved_grant_0,
	WideOr0,
	Equal0,
	Equal11,
	WideOr1,
	m0_write,
	mem_used_7,
	src_data_66,
	out_data_28,
	src_valid,
	src12_valid,
	m0_write1,
	out_data_42,
	out_data_29,
	out_data_31,
	out_data_30,
	out_data_33,
	out_data_32,
	out_data_35,
	out_data_34,
	out_data_37,
	out_data_36,
	out_data_39,
	out_data_38,
	out_data_41,
	out_data_40,
	out_data_19,
	out_data_20,
	out_data_21,
	out_data_22,
	out_data_23,
	out_data_24,
	out_data_25,
	out_data_26,
	out_data_27,
	comb,
	comb1,
	rd_data_0,
	rd_data_1,
	rd_data_2,
	rd_data_3,
	rd_data_4,
	rd_data_5,
	rd_data_6,
	rd_data_7,
	rd_data_8,
	rd_data_9,
	rd_data_10,
	rd_data_11,
	rd_data_12,
	rd_data_13,
	rd_data_14,
	rd_data_15,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	f_select)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	f_pop;
output 	entries_1;
output 	entries_0;
output 	Equal1;
output 	rd_data_27;
output 	rd_data_42;
output 	rd_data_41;
output 	rd_data_28;
output 	rd_data_30;
output 	rd_data_29;
output 	rd_data_32;
output 	rd_data_31;
output 	rd_data_34;
output 	rd_data_33;
output 	rd_data_36;
output 	rd_data_35;
output 	rd_data_38;
output 	rd_data_37;
output 	rd_data_40;
output 	rd_data_39;
input 	Selector41;
output 	rd_data_18;
output 	rd_data_19;
output 	rd_data_20;
output 	rd_data_21;
output 	rd_data_22;
output 	rd_data_23;
output 	rd_data_24;
output 	rd_data_25;
output 	rd_data_26;
output 	rd_data_16;
output 	rd_data_17;
input 	saved_grant_0;
input 	WideOr0;
output 	Equal0;
input 	Equal11;
input 	WideOr1;
input 	m0_write;
input 	mem_used_7;
input 	src_data_66;
input 	out_data_28;
input 	src_valid;
input 	src12_valid;
input 	m0_write1;
input 	out_data_42;
input 	out_data_29;
input 	out_data_31;
input 	out_data_30;
input 	out_data_33;
input 	out_data_32;
input 	out_data_35;
input 	out_data_34;
input 	out_data_37;
input 	out_data_36;
input 	out_data_39;
input 	out_data_38;
input 	out_data_41;
input 	out_data_40;
input 	out_data_19;
input 	out_data_20;
input 	out_data_21;
input 	out_data_22;
input 	out_data_23;
input 	out_data_24;
input 	out_data_25;
input 	out_data_26;
input 	out_data_27;
input 	comb;
input 	comb1;
output 	rd_data_0;
output 	rd_data_1;
output 	rd_data_2;
output 	rd_data_3;
output 	rd_data_4;
output 	rd_data_5;
output 	rd_data_6;
output 	rd_data_7;
output 	rd_data_8;
output 	rd_data_9;
output 	rd_data_10;
output 	rd_data_11;
output 	rd_data_12;
output 	rd_data_13;
output 	rd_data_14;
output 	rd_data_15;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
input 	out_data_5;
input 	out_data_6;
input 	out_data_7;
input 	out_data_8;
input 	out_data_9;
input 	out_data_10;
input 	out_data_11;
input 	out_data_12;
input 	out_data_13;
input 	out_data_14;
input 	out_data_15;
input 	f_select;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always2~0_combout ;
wire \always2~1_combout ;
wire \entries[1]~0_combout ;
wire \entries[0]~1_combout ;
wire \always2~2_combout ;
wire \always2~3_combout ;
wire \wr_address~0_combout ;
wire \wr_address~q ;
wire \entry_1[42]~3_combout ;
wire \entry_1[42]~2_combout ;
wire \entry_1[27]~q ;
wire \entry_0[42]~3_combout ;
wire \entry_0[42]~2_combout ;
wire \entry_0[27]~q ;
wire \rd_address~0_combout ;
wire \rd_address~q ;
wire \entry_1[42]~q ;
wire \entry_0[42]~q ;
wire \entry_1[41]~q ;
wire \entry_0[41]~q ;
wire \entry_1[28]~q ;
wire \entry_0[28]~q ;
wire \entry_1[30]~q ;
wire \entry_0[30]~q ;
wire \entry_1[29]~q ;
wire \entry_0[29]~q ;
wire \entry_1[32]~q ;
wire \entry_0[32]~q ;
wire \entry_1[31]~q ;
wire \entry_0[31]~q ;
wire \entry_1[34]~q ;
wire \entry_0[34]~q ;
wire \entry_1[33]~q ;
wire \entry_0[33]~q ;
wire \entry_1[36]~q ;
wire \entry_0[36]~q ;
wire \entry_1[35]~q ;
wire \entry_0[35]~q ;
wire \entry_1[38]~q ;
wire \entry_0[38]~q ;
wire \entry_1[37]~q ;
wire \entry_0[37]~q ;
wire \entry_1[40]~q ;
wire \entry_0[40]~q ;
wire \entry_1[39]~q ;
wire \entry_0[39]~q ;
wire \entry_1[18]~q ;
wire \entry_0[18]~q ;
wire \entry_1[19]~q ;
wire \entry_0[19]~q ;
wire \entry_1[20]~q ;
wire \entry_0[20]~q ;
wire \entry_1[21]~q ;
wire \entry_0[21]~q ;
wire \entry_1[22]~q ;
wire \entry_0[22]~q ;
wire \entry_1[23]~q ;
wire \entry_0[23]~q ;
wire \entry_1[24]~q ;
wire \entry_0[24]~q ;
wire \entry_1[25]~q ;
wire \entry_0[25]~q ;
wire \entry_1[26]~q ;
wire \entry_0[26]~q ;
wire \entry_1[16]~q ;
wire \entry_0[16]~q ;
wire \entry_1[17]~q ;
wire \entry_0[17]~q ;
wire \entry_1[0]~q ;
wire \entry_0[0]~q ;
wire \entry_1[1]~q ;
wire \entry_0[1]~q ;
wire \entry_1[2]~q ;
wire \entry_0[2]~q ;
wire \entry_1[3]~q ;
wire \entry_0[3]~q ;
wire \entry_1[4]~q ;
wire \entry_0[4]~q ;
wire \entry_1[5]~q ;
wire \entry_0[5]~q ;
wire \entry_1[6]~q ;
wire \entry_0[6]~q ;
wire \entry_1[7]~q ;
wire \entry_0[7]~q ;
wire \entry_1[8]~q ;
wire \entry_0[8]~q ;
wire \entry_1[9]~q ;
wire \entry_0[9]~q ;
wire \entry_1[10]~q ;
wire \entry_0[10]~q ;
wire \entry_1[11]~q ;
wire \entry_0[11]~q ;
wire \entry_1[12]~q ;
wire \entry_0[12]~q ;
wire \entry_1[13]~q ;
wire \entry_0[13]~q ;
wire \entry_1[14]~q ;
wire \entry_0[14]~q ;
wire \entry_1[15]~q ;
wire \entry_0[15]~q ;


dffeas \entries[1] (
	.clk(clk),
	.d(\entries[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(entries_1),
	.prn(vcc));
defparam \entries[1] .is_wysiwyg = "true";
defparam \entries[1] .power_up = "low";

dffeas \entries[0] (
	.clk(clk),
	.d(\entries[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(entries_0),
	.prn(vcc));
defparam \entries[0] .is_wysiwyg = "true";
defparam \entries[0] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEEEE;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[27]~0 (
	.dataa(\entry_1[27]~q ),
	.datab(\entry_0[27]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_27),
	.cout());
defparam \rd_data[27]~0 .lut_mask = 16'hAACC;
defparam \rd_data[27]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[42]~1 (
	.dataa(\entry_1[42]~q ),
	.datab(\entry_0[42]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_42),
	.cout());
defparam \rd_data[42]~1 .lut_mask = 16'hAACC;
defparam \rd_data[42]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[41]~2 (
	.dataa(\entry_1[41]~q ),
	.datab(\entry_0[41]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_41),
	.cout());
defparam \rd_data[41]~2 .lut_mask = 16'hAACC;
defparam \rd_data[41]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[28]~3 (
	.dataa(\entry_1[28]~q ),
	.datab(\entry_0[28]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_28),
	.cout());
defparam \rd_data[28]~3 .lut_mask = 16'hAACC;
defparam \rd_data[28]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[30]~4 (
	.dataa(\entry_1[30]~q ),
	.datab(\entry_0[30]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_30),
	.cout());
defparam \rd_data[30]~4 .lut_mask = 16'hAACC;
defparam \rd_data[30]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[29]~5 (
	.dataa(\entry_1[29]~q ),
	.datab(\entry_0[29]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_29),
	.cout());
defparam \rd_data[29]~5 .lut_mask = 16'hAACC;
defparam \rd_data[29]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[32]~6 (
	.dataa(\entry_1[32]~q ),
	.datab(\entry_0[32]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_32),
	.cout());
defparam \rd_data[32]~6 .lut_mask = 16'hAACC;
defparam \rd_data[32]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[31]~7 (
	.dataa(\entry_1[31]~q ),
	.datab(\entry_0[31]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_31),
	.cout());
defparam \rd_data[31]~7 .lut_mask = 16'hAACC;
defparam \rd_data[31]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[34]~8 (
	.dataa(\entry_1[34]~q ),
	.datab(\entry_0[34]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_34),
	.cout());
defparam \rd_data[34]~8 .lut_mask = 16'hAACC;
defparam \rd_data[34]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[33]~9 (
	.dataa(\entry_1[33]~q ),
	.datab(\entry_0[33]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_33),
	.cout());
defparam \rd_data[33]~9 .lut_mask = 16'hAACC;
defparam \rd_data[33]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[36]~10 (
	.dataa(\entry_1[36]~q ),
	.datab(\entry_0[36]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_36),
	.cout());
defparam \rd_data[36]~10 .lut_mask = 16'hAACC;
defparam \rd_data[36]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[35]~11 (
	.dataa(\entry_1[35]~q ),
	.datab(\entry_0[35]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_35),
	.cout());
defparam \rd_data[35]~11 .lut_mask = 16'hAACC;
defparam \rd_data[35]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[38]~12 (
	.dataa(\entry_1[38]~q ),
	.datab(\entry_0[38]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_38),
	.cout());
defparam \rd_data[38]~12 .lut_mask = 16'hAACC;
defparam \rd_data[38]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[37]~13 (
	.dataa(\entry_1[37]~q ),
	.datab(\entry_0[37]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_37),
	.cout());
defparam \rd_data[37]~13 .lut_mask = 16'hAACC;
defparam \rd_data[37]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[40]~14 (
	.dataa(\entry_1[40]~q ),
	.datab(\entry_0[40]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_40),
	.cout());
defparam \rd_data[40]~14 .lut_mask = 16'hAACC;
defparam \rd_data[40]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[39]~15 (
	.dataa(\entry_1[39]~q ),
	.datab(\entry_0[39]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_39),
	.cout());
defparam \rd_data[39]~15 .lut_mask = 16'hAACC;
defparam \rd_data[39]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[18]~16 (
	.dataa(\entry_1[18]~q ),
	.datab(\entry_0[18]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_18),
	.cout());
defparam \rd_data[18]~16 .lut_mask = 16'hAACC;
defparam \rd_data[18]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[19]~17 (
	.dataa(\entry_1[19]~q ),
	.datab(\entry_0[19]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_19),
	.cout());
defparam \rd_data[19]~17 .lut_mask = 16'hAACC;
defparam \rd_data[19]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[20]~18 (
	.dataa(\entry_1[20]~q ),
	.datab(\entry_0[20]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_20),
	.cout());
defparam \rd_data[20]~18 .lut_mask = 16'hAACC;
defparam \rd_data[20]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[21]~19 (
	.dataa(\entry_1[21]~q ),
	.datab(\entry_0[21]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_21),
	.cout());
defparam \rd_data[21]~19 .lut_mask = 16'hAACC;
defparam \rd_data[21]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[22]~20 (
	.dataa(\entry_1[22]~q ),
	.datab(\entry_0[22]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_22),
	.cout());
defparam \rd_data[22]~20 .lut_mask = 16'hAACC;
defparam \rd_data[22]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[23]~21 (
	.dataa(\entry_1[23]~q ),
	.datab(\entry_0[23]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_23),
	.cout());
defparam \rd_data[23]~21 .lut_mask = 16'hAACC;
defparam \rd_data[23]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[24]~22 (
	.dataa(\entry_1[24]~q ),
	.datab(\entry_0[24]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_24),
	.cout());
defparam \rd_data[24]~22 .lut_mask = 16'hAACC;
defparam \rd_data[24]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[25]~23 (
	.dataa(\entry_1[25]~q ),
	.datab(\entry_0[25]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_25),
	.cout());
defparam \rd_data[25]~23 .lut_mask = 16'hAACC;
defparam \rd_data[25]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[26]~24 (
	.dataa(\entry_1[26]~q ),
	.datab(\entry_0[26]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_26),
	.cout());
defparam \rd_data[26]~24 .lut_mask = 16'hAACC;
defparam \rd_data[26]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[16]~25 (
	.dataa(\entry_1[16]~q ),
	.datab(\entry_0[16]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_16),
	.cout());
defparam \rd_data[16]~25 .lut_mask = 16'hAACC;
defparam \rd_data[16]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[17]~26 (
	.dataa(\entry_1[17]~q ),
	.datab(\entry_0[17]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_17),
	.cout());
defparam \rd_data[17]~26 .lut_mask = 16'hAACC;
defparam \rd_data[17]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(entries_1),
	.datab(gnd),
	.datac(gnd),
	.datad(entries_0),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hAAFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[0]~27 (
	.dataa(\entry_1[0]~q ),
	.datab(\entry_0[0]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_0),
	.cout());
defparam \rd_data[0]~27 .lut_mask = 16'hAACC;
defparam \rd_data[0]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[1]~28 (
	.dataa(\entry_1[1]~q ),
	.datab(\entry_0[1]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_1),
	.cout());
defparam \rd_data[1]~28 .lut_mask = 16'hAACC;
defparam \rd_data[1]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[2]~29 (
	.dataa(\entry_1[2]~q ),
	.datab(\entry_0[2]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_2),
	.cout());
defparam \rd_data[2]~29 .lut_mask = 16'hAACC;
defparam \rd_data[2]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[3]~30 (
	.dataa(\entry_1[3]~q ),
	.datab(\entry_0[3]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_3),
	.cout());
defparam \rd_data[3]~30 .lut_mask = 16'hAACC;
defparam \rd_data[3]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[4]~31 (
	.dataa(\entry_1[4]~q ),
	.datab(\entry_0[4]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_4),
	.cout());
defparam \rd_data[4]~31 .lut_mask = 16'hAACC;
defparam \rd_data[4]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[5]~32 (
	.dataa(\entry_1[5]~q ),
	.datab(\entry_0[5]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_5),
	.cout());
defparam \rd_data[5]~32 .lut_mask = 16'hAACC;
defparam \rd_data[5]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[6]~33 (
	.dataa(\entry_1[6]~q ),
	.datab(\entry_0[6]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_6),
	.cout());
defparam \rd_data[6]~33 .lut_mask = 16'hAACC;
defparam \rd_data[6]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[7]~34 (
	.dataa(\entry_1[7]~q ),
	.datab(\entry_0[7]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_7),
	.cout());
defparam \rd_data[7]~34 .lut_mask = 16'hAACC;
defparam \rd_data[7]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[8]~35 (
	.dataa(\entry_1[8]~q ),
	.datab(\entry_0[8]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_8),
	.cout());
defparam \rd_data[8]~35 .lut_mask = 16'hAACC;
defparam \rd_data[8]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[9]~36 (
	.dataa(\entry_1[9]~q ),
	.datab(\entry_0[9]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_9),
	.cout());
defparam \rd_data[9]~36 .lut_mask = 16'hAACC;
defparam \rd_data[9]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[10]~37 (
	.dataa(\entry_1[10]~q ),
	.datab(\entry_0[10]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_10),
	.cout());
defparam \rd_data[10]~37 .lut_mask = 16'hAACC;
defparam \rd_data[10]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[11]~38 (
	.dataa(\entry_1[11]~q ),
	.datab(\entry_0[11]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_11),
	.cout());
defparam \rd_data[11]~38 .lut_mask = 16'hAACC;
defparam \rd_data[11]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[12]~39 (
	.dataa(\entry_1[12]~q ),
	.datab(\entry_0[12]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_12),
	.cout());
defparam \rd_data[12]~39 .lut_mask = 16'hAACC;
defparam \rd_data[12]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[13]~40 (
	.dataa(\entry_1[13]~q ),
	.datab(\entry_0[13]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_13),
	.cout());
defparam \rd_data[13]~40 .lut_mask = 16'hAACC;
defparam \rd_data[13]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[14]~41 (
	.dataa(\entry_1[14]~q ),
	.datab(\entry_0[14]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_14),
	.cout());
defparam \rd_data[14]~41 .lut_mask = 16'hAACC;
defparam \rd_data[14]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[15]~42 (
	.dataa(\entry_1[15]~q ),
	.datab(\entry_0[15]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_15),
	.cout());
defparam \rd_data[15]~42 .lut_mask = 16'hAACC;
defparam \rd_data[15]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(m0_write),
	.datab(mem_used_7),
	.datac(src_data_66),
	.datad(gnd),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hFBFB;
defparam \always2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~1 (
	.dataa(WideOr0),
	.datab(Equal0),
	.datac(WideOr1),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\always2~1_combout ),
	.cout());
defparam \always2~1 .lut_mask = 16'hFFFB;
defparam \always2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \entries[1]~0 (
	.dataa(entries_1),
	.datab(f_select),
	.datac(entries_0),
	.datad(\always2~1_combout ),
	.cin(gnd),
	.combout(\entries[1]~0_combout ),
	.cout());
defparam \entries[1]~0 .lut_mask = 16'h6996;
defparam \entries[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \entries[0]~1 (
	.dataa(entries_0),
	.datab(f_select),
	.datac(\always2~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\entries[0]~1_combout ),
	.cout());
defparam \entries[0]~1 .lut_mask = 16'h9696;
defparam \entries[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~2 (
	.dataa(src_data_66),
	.datab(mem_used_7),
	.datac(src_valid),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(\always2~2_combout ),
	.cout());
defparam \always2~2 .lut_mask = 16'hFFFB;
defparam \always2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~3 (
	.dataa(src_valid),
	.datab(src12_valid),
	.datac(Equal11),
	.datad(\always2~2_combout ),
	.cin(gnd),
	.combout(\always2~3_combout ),
	.cout());
defparam \always2~3 .lut_mask = 16'hFFEF;
defparam \always2~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_address~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\always2~1_combout ),
	.datad(\wr_address~q ),
	.cin(gnd),
	.combout(\wr_address~0_combout ),
	.cout());
defparam \wr_address~0 .lut_mask = 16'h0FF0;
defparam \wr_address~0 .sum_lutc_input = "datac";

dffeas wr_address(
	.clk(clk),
	.d(\wr_address~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_address~q ),
	.prn(vcc));
defparam wr_address.is_wysiwyg = "true";
defparam wr_address.power_up = "low";

cycloneive_lcell_comb \entry_1[42]~3 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\wr_address~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\entry_1[42]~3_combout ),
	.cout());
defparam \entry_1[42]~3 .lut_mask = 16'hFDFD;
defparam \entry_1[42]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \entry_1[42]~2 (
	.dataa(m0_write1),
	.datab(\always2~3_combout ),
	.datac(WideOr0),
	.datad(\entry_1[42]~3_combout ),
	.cin(gnd),
	.combout(\entry_1[42]~2_combout ),
	.cout());
defparam \entry_1[42]~2 .lut_mask = 16'hFFFD;
defparam \entry_1[42]~2 .sum_lutc_input = "datac";

dffeas \entry_1[27] (
	.clk(clk),
	.d(out_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[27]~q ),
	.prn(vcc));
defparam \entry_1[27] .is_wysiwyg = "true";
defparam \entry_1[27] .power_up = "low";

cycloneive_lcell_comb \entry_0[42]~3 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\wr_address~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\entry_0[42]~3_combout ),
	.cout());
defparam \entry_0[42]~3 .lut_mask = 16'hDFDF;
defparam \entry_0[42]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \entry_0[42]~2 (
	.dataa(m0_write1),
	.datab(\always2~3_combout ),
	.datac(WideOr0),
	.datad(\entry_0[42]~3_combout ),
	.cin(gnd),
	.combout(\entry_0[42]~2_combout ),
	.cout());
defparam \entry_0[42]~2 .lut_mask = 16'hFFFD;
defparam \entry_0[42]~2 .sum_lutc_input = "datac";

dffeas \entry_0[27] (
	.clk(clk),
	.d(out_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[27]~q ),
	.prn(vcc));
defparam \entry_0[27] .is_wysiwyg = "true";
defparam \entry_0[27] .power_up = "low";

cycloneive_lcell_comb \rd_address~0 (
	.dataa(gnd),
	.datab(\rd_address~q ),
	.datac(f_pop),
	.datad(Selector41),
	.cin(gnd),
	.combout(\rd_address~0_combout ),
	.cout());
defparam \rd_address~0 .lut_mask = 16'hC33C;
defparam \rd_address~0 .sum_lutc_input = "datac";

dffeas rd_address(
	.clk(clk),
	.d(\rd_address~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_address~q ),
	.prn(vcc));
defparam rd_address.is_wysiwyg = "true";
defparam rd_address.power_up = "low";

dffeas \entry_1[42] (
	.clk(clk),
	.d(m0_write1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[42]~q ),
	.prn(vcc));
defparam \entry_1[42] .is_wysiwyg = "true";
defparam \entry_1[42] .power_up = "low";

dffeas \entry_0[42] (
	.clk(clk),
	.d(m0_write1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[42]~q ),
	.prn(vcc));
defparam \entry_0[42] .is_wysiwyg = "true";
defparam \entry_0[42] .power_up = "low";

dffeas \entry_1[41] (
	.clk(clk),
	.d(out_data_42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[41]~q ),
	.prn(vcc));
defparam \entry_1[41] .is_wysiwyg = "true";
defparam \entry_1[41] .power_up = "low";

dffeas \entry_0[41] (
	.clk(clk),
	.d(out_data_42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[41]~q ),
	.prn(vcc));
defparam \entry_0[41] .is_wysiwyg = "true";
defparam \entry_0[41] .power_up = "low";

dffeas \entry_1[28] (
	.clk(clk),
	.d(out_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[28]~q ),
	.prn(vcc));
defparam \entry_1[28] .is_wysiwyg = "true";
defparam \entry_1[28] .power_up = "low";

dffeas \entry_0[28] (
	.clk(clk),
	.d(out_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[28]~q ),
	.prn(vcc));
defparam \entry_0[28] .is_wysiwyg = "true";
defparam \entry_0[28] .power_up = "low";

dffeas \entry_1[30] (
	.clk(clk),
	.d(out_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[30]~q ),
	.prn(vcc));
defparam \entry_1[30] .is_wysiwyg = "true";
defparam \entry_1[30] .power_up = "low";

dffeas \entry_0[30] (
	.clk(clk),
	.d(out_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[30]~q ),
	.prn(vcc));
defparam \entry_0[30] .is_wysiwyg = "true";
defparam \entry_0[30] .power_up = "low";

dffeas \entry_1[29] (
	.clk(clk),
	.d(out_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[29]~q ),
	.prn(vcc));
defparam \entry_1[29] .is_wysiwyg = "true";
defparam \entry_1[29] .power_up = "low";

dffeas \entry_0[29] (
	.clk(clk),
	.d(out_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[29]~q ),
	.prn(vcc));
defparam \entry_0[29] .is_wysiwyg = "true";
defparam \entry_0[29] .power_up = "low";

dffeas \entry_1[32] (
	.clk(clk),
	.d(out_data_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[32]~q ),
	.prn(vcc));
defparam \entry_1[32] .is_wysiwyg = "true";
defparam \entry_1[32] .power_up = "low";

dffeas \entry_0[32] (
	.clk(clk),
	.d(out_data_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[32]~q ),
	.prn(vcc));
defparam \entry_0[32] .is_wysiwyg = "true";
defparam \entry_0[32] .power_up = "low";

dffeas \entry_1[31] (
	.clk(clk),
	.d(out_data_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[31]~q ),
	.prn(vcc));
defparam \entry_1[31] .is_wysiwyg = "true";
defparam \entry_1[31] .power_up = "low";

dffeas \entry_0[31] (
	.clk(clk),
	.d(out_data_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[31]~q ),
	.prn(vcc));
defparam \entry_0[31] .is_wysiwyg = "true";
defparam \entry_0[31] .power_up = "low";

dffeas \entry_1[34] (
	.clk(clk),
	.d(out_data_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[34]~q ),
	.prn(vcc));
defparam \entry_1[34] .is_wysiwyg = "true";
defparam \entry_1[34] .power_up = "low";

dffeas \entry_0[34] (
	.clk(clk),
	.d(out_data_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[34]~q ),
	.prn(vcc));
defparam \entry_0[34] .is_wysiwyg = "true";
defparam \entry_0[34] .power_up = "low";

dffeas \entry_1[33] (
	.clk(clk),
	.d(out_data_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[33]~q ),
	.prn(vcc));
defparam \entry_1[33] .is_wysiwyg = "true";
defparam \entry_1[33] .power_up = "low";

dffeas \entry_0[33] (
	.clk(clk),
	.d(out_data_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[33]~q ),
	.prn(vcc));
defparam \entry_0[33] .is_wysiwyg = "true";
defparam \entry_0[33] .power_up = "low";

dffeas \entry_1[36] (
	.clk(clk),
	.d(out_data_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[36]~q ),
	.prn(vcc));
defparam \entry_1[36] .is_wysiwyg = "true";
defparam \entry_1[36] .power_up = "low";

dffeas \entry_0[36] (
	.clk(clk),
	.d(out_data_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[36]~q ),
	.prn(vcc));
defparam \entry_0[36] .is_wysiwyg = "true";
defparam \entry_0[36] .power_up = "low";

dffeas \entry_1[35] (
	.clk(clk),
	.d(out_data_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[35]~q ),
	.prn(vcc));
defparam \entry_1[35] .is_wysiwyg = "true";
defparam \entry_1[35] .power_up = "low";

dffeas \entry_0[35] (
	.clk(clk),
	.d(out_data_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[35]~q ),
	.prn(vcc));
defparam \entry_0[35] .is_wysiwyg = "true";
defparam \entry_0[35] .power_up = "low";

dffeas \entry_1[38] (
	.clk(clk),
	.d(out_data_39),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[38]~q ),
	.prn(vcc));
defparam \entry_1[38] .is_wysiwyg = "true";
defparam \entry_1[38] .power_up = "low";

dffeas \entry_0[38] (
	.clk(clk),
	.d(out_data_39),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[38]~q ),
	.prn(vcc));
defparam \entry_0[38] .is_wysiwyg = "true";
defparam \entry_0[38] .power_up = "low";

dffeas \entry_1[37] (
	.clk(clk),
	.d(out_data_38),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[37]~q ),
	.prn(vcc));
defparam \entry_1[37] .is_wysiwyg = "true";
defparam \entry_1[37] .power_up = "low";

dffeas \entry_0[37] (
	.clk(clk),
	.d(out_data_38),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[37]~q ),
	.prn(vcc));
defparam \entry_0[37] .is_wysiwyg = "true";
defparam \entry_0[37] .power_up = "low";

dffeas \entry_1[40] (
	.clk(clk),
	.d(out_data_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[40]~q ),
	.prn(vcc));
defparam \entry_1[40] .is_wysiwyg = "true";
defparam \entry_1[40] .power_up = "low";

dffeas \entry_0[40] (
	.clk(clk),
	.d(out_data_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[40]~q ),
	.prn(vcc));
defparam \entry_0[40] .is_wysiwyg = "true";
defparam \entry_0[40] .power_up = "low";

dffeas \entry_1[39] (
	.clk(clk),
	.d(out_data_40),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[39]~q ),
	.prn(vcc));
defparam \entry_1[39] .is_wysiwyg = "true";
defparam \entry_1[39] .power_up = "low";

dffeas \entry_0[39] (
	.clk(clk),
	.d(out_data_40),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[39]~q ),
	.prn(vcc));
defparam \entry_0[39] .is_wysiwyg = "true";
defparam \entry_0[39] .power_up = "low";

dffeas \entry_1[18] (
	.clk(clk),
	.d(out_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[18]~q ),
	.prn(vcc));
defparam \entry_1[18] .is_wysiwyg = "true";
defparam \entry_1[18] .power_up = "low";

dffeas \entry_0[18] (
	.clk(clk),
	.d(out_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[18]~q ),
	.prn(vcc));
defparam \entry_0[18] .is_wysiwyg = "true";
defparam \entry_0[18] .power_up = "low";

dffeas \entry_1[19] (
	.clk(clk),
	.d(out_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[19]~q ),
	.prn(vcc));
defparam \entry_1[19] .is_wysiwyg = "true";
defparam \entry_1[19] .power_up = "low";

dffeas \entry_0[19] (
	.clk(clk),
	.d(out_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[19]~q ),
	.prn(vcc));
defparam \entry_0[19] .is_wysiwyg = "true";
defparam \entry_0[19] .power_up = "low";

dffeas \entry_1[20] (
	.clk(clk),
	.d(out_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[20]~q ),
	.prn(vcc));
defparam \entry_1[20] .is_wysiwyg = "true";
defparam \entry_1[20] .power_up = "low";

dffeas \entry_0[20] (
	.clk(clk),
	.d(out_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[20]~q ),
	.prn(vcc));
defparam \entry_0[20] .is_wysiwyg = "true";
defparam \entry_0[20] .power_up = "low";

dffeas \entry_1[21] (
	.clk(clk),
	.d(out_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[21]~q ),
	.prn(vcc));
defparam \entry_1[21] .is_wysiwyg = "true";
defparam \entry_1[21] .power_up = "low";

dffeas \entry_0[21] (
	.clk(clk),
	.d(out_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[21]~q ),
	.prn(vcc));
defparam \entry_0[21] .is_wysiwyg = "true";
defparam \entry_0[21] .power_up = "low";

dffeas \entry_1[22] (
	.clk(clk),
	.d(out_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[22]~q ),
	.prn(vcc));
defparam \entry_1[22] .is_wysiwyg = "true";
defparam \entry_1[22] .power_up = "low";

dffeas \entry_0[22] (
	.clk(clk),
	.d(out_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[22]~q ),
	.prn(vcc));
defparam \entry_0[22] .is_wysiwyg = "true";
defparam \entry_0[22] .power_up = "low";

dffeas \entry_1[23] (
	.clk(clk),
	.d(out_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[23]~q ),
	.prn(vcc));
defparam \entry_1[23] .is_wysiwyg = "true";
defparam \entry_1[23] .power_up = "low";

dffeas \entry_0[23] (
	.clk(clk),
	.d(out_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[23]~q ),
	.prn(vcc));
defparam \entry_0[23] .is_wysiwyg = "true";
defparam \entry_0[23] .power_up = "low";

dffeas \entry_1[24] (
	.clk(clk),
	.d(out_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[24]~q ),
	.prn(vcc));
defparam \entry_1[24] .is_wysiwyg = "true";
defparam \entry_1[24] .power_up = "low";

dffeas \entry_0[24] (
	.clk(clk),
	.d(out_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[24]~q ),
	.prn(vcc));
defparam \entry_0[24] .is_wysiwyg = "true";
defparam \entry_0[24] .power_up = "low";

dffeas \entry_1[25] (
	.clk(clk),
	.d(out_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[25]~q ),
	.prn(vcc));
defparam \entry_1[25] .is_wysiwyg = "true";
defparam \entry_1[25] .power_up = "low";

dffeas \entry_0[25] (
	.clk(clk),
	.d(out_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[25]~q ),
	.prn(vcc));
defparam \entry_0[25] .is_wysiwyg = "true";
defparam \entry_0[25] .power_up = "low";

dffeas \entry_1[26] (
	.clk(clk),
	.d(out_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[26]~q ),
	.prn(vcc));
defparam \entry_1[26] .is_wysiwyg = "true";
defparam \entry_1[26] .power_up = "low";

dffeas \entry_0[26] (
	.clk(clk),
	.d(out_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[26]~q ),
	.prn(vcc));
defparam \entry_0[26] .is_wysiwyg = "true";
defparam \entry_0[26] .power_up = "low";

dffeas \entry_1[16] (
	.clk(clk),
	.d(comb),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[16]~q ),
	.prn(vcc));
defparam \entry_1[16] .is_wysiwyg = "true";
defparam \entry_1[16] .power_up = "low";

dffeas \entry_0[16] (
	.clk(clk),
	.d(comb),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[16]~q ),
	.prn(vcc));
defparam \entry_0[16] .is_wysiwyg = "true";
defparam \entry_0[16] .power_up = "low";

dffeas \entry_1[17] (
	.clk(clk),
	.d(comb1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[17]~q ),
	.prn(vcc));
defparam \entry_1[17] .is_wysiwyg = "true";
defparam \entry_1[17] .power_up = "low";

dffeas \entry_0[17] (
	.clk(clk),
	.d(comb1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[17]~q ),
	.prn(vcc));
defparam \entry_0[17] .is_wysiwyg = "true";
defparam \entry_0[17] .power_up = "low";

dffeas \entry_1[0] (
	.clk(clk),
	.d(out_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[0]~q ),
	.prn(vcc));
defparam \entry_1[0] .is_wysiwyg = "true";
defparam \entry_1[0] .power_up = "low";

dffeas \entry_0[0] (
	.clk(clk),
	.d(out_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[0]~q ),
	.prn(vcc));
defparam \entry_0[0] .is_wysiwyg = "true";
defparam \entry_0[0] .power_up = "low";

dffeas \entry_1[1] (
	.clk(clk),
	.d(out_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[1]~q ),
	.prn(vcc));
defparam \entry_1[1] .is_wysiwyg = "true";
defparam \entry_1[1] .power_up = "low";

dffeas \entry_0[1] (
	.clk(clk),
	.d(out_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[1]~q ),
	.prn(vcc));
defparam \entry_0[1] .is_wysiwyg = "true";
defparam \entry_0[1] .power_up = "low";

dffeas \entry_1[2] (
	.clk(clk),
	.d(out_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[2]~q ),
	.prn(vcc));
defparam \entry_1[2] .is_wysiwyg = "true";
defparam \entry_1[2] .power_up = "low";

dffeas \entry_0[2] (
	.clk(clk),
	.d(out_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[2]~q ),
	.prn(vcc));
defparam \entry_0[2] .is_wysiwyg = "true";
defparam \entry_0[2] .power_up = "low";

dffeas \entry_1[3] (
	.clk(clk),
	.d(out_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[3]~q ),
	.prn(vcc));
defparam \entry_1[3] .is_wysiwyg = "true";
defparam \entry_1[3] .power_up = "low";

dffeas \entry_0[3] (
	.clk(clk),
	.d(out_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[3]~q ),
	.prn(vcc));
defparam \entry_0[3] .is_wysiwyg = "true";
defparam \entry_0[3] .power_up = "low";

dffeas \entry_1[4] (
	.clk(clk),
	.d(out_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[4]~q ),
	.prn(vcc));
defparam \entry_1[4] .is_wysiwyg = "true";
defparam \entry_1[4] .power_up = "low";

dffeas \entry_0[4] (
	.clk(clk),
	.d(out_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[4]~q ),
	.prn(vcc));
defparam \entry_0[4] .is_wysiwyg = "true";
defparam \entry_0[4] .power_up = "low";

dffeas \entry_1[5] (
	.clk(clk),
	.d(out_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[5]~q ),
	.prn(vcc));
defparam \entry_1[5] .is_wysiwyg = "true";
defparam \entry_1[5] .power_up = "low";

dffeas \entry_0[5] (
	.clk(clk),
	.d(out_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[5]~q ),
	.prn(vcc));
defparam \entry_0[5] .is_wysiwyg = "true";
defparam \entry_0[5] .power_up = "low";

dffeas \entry_1[6] (
	.clk(clk),
	.d(out_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[6]~q ),
	.prn(vcc));
defparam \entry_1[6] .is_wysiwyg = "true";
defparam \entry_1[6] .power_up = "low";

dffeas \entry_0[6] (
	.clk(clk),
	.d(out_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[6]~q ),
	.prn(vcc));
defparam \entry_0[6] .is_wysiwyg = "true";
defparam \entry_0[6] .power_up = "low";

dffeas \entry_1[7] (
	.clk(clk),
	.d(out_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[7]~q ),
	.prn(vcc));
defparam \entry_1[7] .is_wysiwyg = "true";
defparam \entry_1[7] .power_up = "low";

dffeas \entry_0[7] (
	.clk(clk),
	.d(out_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[7]~q ),
	.prn(vcc));
defparam \entry_0[7] .is_wysiwyg = "true";
defparam \entry_0[7] .power_up = "low";

dffeas \entry_1[8] (
	.clk(clk),
	.d(out_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[8]~q ),
	.prn(vcc));
defparam \entry_1[8] .is_wysiwyg = "true";
defparam \entry_1[8] .power_up = "low";

dffeas \entry_0[8] (
	.clk(clk),
	.d(out_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[8]~q ),
	.prn(vcc));
defparam \entry_0[8] .is_wysiwyg = "true";
defparam \entry_0[8] .power_up = "low";

dffeas \entry_1[9] (
	.clk(clk),
	.d(out_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[9]~q ),
	.prn(vcc));
defparam \entry_1[9] .is_wysiwyg = "true";
defparam \entry_1[9] .power_up = "low";

dffeas \entry_0[9] (
	.clk(clk),
	.d(out_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[9]~q ),
	.prn(vcc));
defparam \entry_0[9] .is_wysiwyg = "true";
defparam \entry_0[9] .power_up = "low";

dffeas \entry_1[10] (
	.clk(clk),
	.d(out_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[10]~q ),
	.prn(vcc));
defparam \entry_1[10] .is_wysiwyg = "true";
defparam \entry_1[10] .power_up = "low";

dffeas \entry_0[10] (
	.clk(clk),
	.d(out_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[10]~q ),
	.prn(vcc));
defparam \entry_0[10] .is_wysiwyg = "true";
defparam \entry_0[10] .power_up = "low";

dffeas \entry_1[11] (
	.clk(clk),
	.d(out_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[11]~q ),
	.prn(vcc));
defparam \entry_1[11] .is_wysiwyg = "true";
defparam \entry_1[11] .power_up = "low";

dffeas \entry_0[11] (
	.clk(clk),
	.d(out_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[11]~q ),
	.prn(vcc));
defparam \entry_0[11] .is_wysiwyg = "true";
defparam \entry_0[11] .power_up = "low";

dffeas \entry_1[12] (
	.clk(clk),
	.d(out_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[12]~q ),
	.prn(vcc));
defparam \entry_1[12] .is_wysiwyg = "true";
defparam \entry_1[12] .power_up = "low";

dffeas \entry_0[12] (
	.clk(clk),
	.d(out_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[12]~q ),
	.prn(vcc));
defparam \entry_0[12] .is_wysiwyg = "true";
defparam \entry_0[12] .power_up = "low";

dffeas \entry_1[13] (
	.clk(clk),
	.d(out_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[13]~q ),
	.prn(vcc));
defparam \entry_1[13] .is_wysiwyg = "true";
defparam \entry_1[13] .power_up = "low";

dffeas \entry_0[13] (
	.clk(clk),
	.d(out_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[13]~q ),
	.prn(vcc));
defparam \entry_0[13] .is_wysiwyg = "true";
defparam \entry_0[13] .power_up = "low";

dffeas \entry_1[14] (
	.clk(clk),
	.d(out_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[14]~q ),
	.prn(vcc));
defparam \entry_1[14] .is_wysiwyg = "true";
defparam \entry_1[14] .power_up = "low";

dffeas \entry_0[14] (
	.clk(clk),
	.d(out_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[14]~q ),
	.prn(vcc));
defparam \entry_0[14] .is_wysiwyg = "true";
defparam \entry_0[14] .power_up = "low";

dffeas \entry_1[15] (
	.clk(clk),
	.d(out_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[42]~2_combout ),
	.q(\entry_1[15]~q ),
	.prn(vcc));
defparam \entry_1[15] .is_wysiwyg = "true";
defparam \entry_1[15] .power_up = "low";

dffeas \entry_0[15] (
	.clk(clk),
	.d(out_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[42]~2_combout ),
	.q(\entry_0[15]~q ),
	.prn(vcc));
defparam \entry_0[15] .is_wysiwyg = "true";
defparam \entry_0[15] .power_up = "low";

endmodule

module niosII_niosII_sys_pll (
	wire_pll7_clk_0,
	wire_pll7_clk_1,
	out_data_buffer_0,
	out_data_toggle_flopped,
	dreg_0,
	mem_used_1,
	wire_pfdena_reg_ena,
	out_data_buffer_65,
	out_data_buffer_38,
	out_data_buffer_39,
	reset,
	out_data_buffer_66,
	readdata_0,
	readdata_1,
	out_data_buffer_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	wire_pll7_clk_0;
output 	wire_pll7_clk_1;
input 	out_data_buffer_0;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	mem_used_1;
output 	wire_pfdena_reg_ena;
input 	out_data_buffer_65;
input 	out_data_buffer_38;
input 	out_data_buffer_39;
input 	reset;
input 	out_data_buffer_66;
output 	readdata_0;
output 	readdata_1;
input 	out_data_buffer_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \stdsync2|dffpipe3|dffe6a[0]~q ;
wire \sd1|locked~combout ;
wire \readdata[0]~0_combout ;
wire \wire_pfdena_reg_ena~1_combout ;
wire \w_reset~combout ;
wire \prev_reset~q ;
wire \pfdena_reg~0_combout ;
wire \pfdena_reg~q ;


niosII_niosII_sys_pll_altpll_8ra2 sd1(
	.clk({clk_unconnected_wire_4,clk_unconnected_wire_3,clk_unconnected_wire_2,wire_pll7_clk_1,wire_pll7_clk_0}),
	.areset(\prev_reset~q ),
	.locked1(\sd1|locked~combout ),
	.inclk({gnd,clk_clk}));

niosII_niosII_sys_pll_stdsync_sv6 stdsync2(
	.altera_reset_synchronizer_int_chain_out(reset),
	.dffe6a_0(\stdsync2|dffpipe3|dffe6a[0]~q ),
	.locked(\sd1|locked~combout ),
	.clk_clk(clk_clk));

cycloneive_lcell_comb \wire_pfdena_reg_ena~0 (
	.dataa(gnd),
	.datab(out_data_toggle_flopped),
	.datac(dreg_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(wire_pfdena_reg_ena),
	.cout());
defparam \wire_pfdena_reg_ena~0 .lut_mask = 16'h3CFF;
defparam \wire_pfdena_reg_ena~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0]~1 (
	.dataa(\readdata[0]~0_combout ),
	.datab(\prev_reset~q ),
	.datac(\stdsync2|dffpipe3|dffe6a[0]~q ),
	.datad(out_data_buffer_38),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0]~1 .lut_mask = 16'hFAFC;
defparam \readdata[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1]~2 (
	.dataa(\readdata[0]~0_combout ),
	.datab(gnd),
	.datac(out_data_buffer_38),
	.datad(\pfdena_reg~q ),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1]~2 .lut_mask = 16'hAFFF;
defparam \readdata[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0]~0 (
	.dataa(wire_pfdena_reg_ena),
	.datab(out_data_buffer_66),
	.datac(gnd),
	.datad(out_data_buffer_39),
	.cin(gnd),
	.combout(\readdata[0]~0_combout ),
	.cout());
defparam \readdata[0]~0 .lut_mask = 16'hEEFF;
defparam \readdata[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wire_pfdena_reg_ena~1 (
	.dataa(wire_pfdena_reg_ena),
	.datab(out_data_buffer_65),
	.datac(out_data_buffer_38),
	.datad(out_data_buffer_39),
	.cin(gnd),
	.combout(\wire_pfdena_reg_ena~1_combout ),
	.cout());
defparam \wire_pfdena_reg_ena~1 .lut_mask = 16'hFEFF;
defparam \wire_pfdena_reg_ena~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb w_reset(
	.dataa(out_data_buffer_0),
	.datab(\wire_pfdena_reg_ena~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\w_reset~combout ),
	.cout());
defparam w_reset.lut_mask = 16'hEEEE;
defparam w_reset.sum_lutc_input = "datac";

dffeas prev_reset(
	.clk(clk_clk),
	.d(\w_reset~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\prev_reset~q ),
	.prn(vcc));
defparam prev_reset.is_wysiwyg = "true";
defparam prev_reset.power_up = "low";

cycloneive_lcell_comb \pfdena_reg~0 (
	.dataa(out_data_buffer_1),
	.datab(\wire_pfdena_reg_ena~1_combout ),
	.datac(gnd),
	.datad(\pfdena_reg~q ),
	.cin(gnd),
	.combout(\pfdena_reg~0_combout ),
	.cout());
defparam \pfdena_reg~0 .lut_mask = 16'hDD11;
defparam \pfdena_reg~0 .sum_lutc_input = "datac";

dffeas pfdena_reg(
	.clk(clk_clk),
	.d(\pfdena_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pfdena_reg~q ),
	.prn(vcc));
defparam pfdena_reg.is_wysiwyg = "true";
defparam pfdena_reg.power_up = "low";

endmodule

module niosII_niosII_sys_pll_altpll_8ra2 (
	clk,
	areset,
	locked1,
	inclk)/* synthesis synthesis_greybox=1 */;
output 	[4:0] clk;
input 	areset;
output 	locked1;
input 	[1:0] inclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wire_pll7_clk[2] ;
wire \wire_pll7_clk[3] ;
wire \wire_pll7_clk[4] ;
wire wire_pll7_locked;
wire wire_pll7_fbout;
wire \pll_lock_sync~q ;

wire [4:0] pll7_CLK_bus;

assign clk[0] = pll7_CLK_bus[0];
assign clk[1] = pll7_CLK_bus[1];
assign \wire_pll7_clk[2]  = pll7_CLK_bus[2];
assign \wire_pll7_clk[3]  = pll7_CLK_bus[3];
assign \wire_pll7_clk[4]  = pll7_CLK_bus[4];

cycloneive_pll pll7(
	.areset(areset),
	.pfdena(vcc),
	.fbin(wire_pll7_fbout),
	.phaseupdown(gnd),
	.phasestep(gnd),
	.scandata(gnd),
	.scanclk(gnd),
	.scanclkena(vcc),
	.configupdate(gnd),
	.clkswitch(gnd),
	.inclk({gnd,inclk[0]}),
	.phasecounterselect(3'b000),
	.phasedone(),
	.scandataout(),
	.scandone(),
	.activeclock(),
	.locked(wire_pll7_locked),
	.vcooverrange(),
	.vcounderrange(),
	.fbout(wire_pll7_fbout),
	.clk(pll7_CLK_bus),
	.clkbad());
defparam pll7.auto_settings = "false";
defparam pll7.bandwidth_type = "auto";
defparam pll7.c0_high = 5;
defparam pll7.c0_initial = 2;
defparam pll7.c0_low = 4;
defparam pll7.c0_mode = "odd";
defparam pll7.c0_ph = 4;
defparam pll7.c1_high = 5;
defparam pll7.c1_initial = 1;
defparam pll7.c1_low = 4;
defparam pll7.c1_mode = "odd";
defparam pll7.c1_ph = 0;
defparam pll7.c1_use_casc_in = "off";
defparam pll7.c2_high = 1;
defparam pll7.c2_initial = 1;
defparam pll7.c2_low = 1;
defparam pll7.c2_mode = "bypass";
defparam pll7.c2_ph = 0;
defparam pll7.c2_use_casc_in = "off";
defparam pll7.c3_high = 1;
defparam pll7.c3_initial = 1;
defparam pll7.c3_low = 1;
defparam pll7.c3_mode = "bypass";
defparam pll7.c3_ph = 0;
defparam pll7.c3_use_casc_in = "off";
defparam pll7.c4_high = 1;
defparam pll7.c4_initial = 1;
defparam pll7.c4_low = 1;
defparam pll7.c4_mode = "bypass";
defparam pll7.c4_ph = 0;
defparam pll7.c4_use_casc_in = "off";
defparam pll7.charge_pump_current_bits = 2;
defparam pll7.clk0_counter = "c0";
defparam pll7.clk0_divide_by = 1;
defparam pll7.clk0_duty_cycle = 50;
defparam pll7.clk0_multiply_by = 2;
defparam pll7.clk0_phase_shift = "0";
defparam pll7.clk1_counter = "c1";
defparam pll7.clk1_divide_by = 1;
defparam pll7.clk1_duty_cycle = 50;
defparam pll7.clk1_multiply_by = 2;
defparam pll7.clk1_phase_shift = "-1667";
defparam pll7.clk2_counter = "unused";
defparam pll7.clk2_divide_by = 0;
defparam pll7.clk2_duty_cycle = 50;
defparam pll7.clk2_multiply_by = 0;
defparam pll7.clk2_phase_shift = "0";
defparam pll7.clk3_counter = "unused";
defparam pll7.clk3_divide_by = 0;
defparam pll7.clk3_duty_cycle = 50;
defparam pll7.clk3_multiply_by = 0;
defparam pll7.clk3_phase_shift = "0";
defparam pll7.clk4_counter = "unused";
defparam pll7.clk4_divide_by = 0;
defparam pll7.clk4_duty_cycle = 50;
defparam pll7.clk4_multiply_by = 0;
defparam pll7.clk4_phase_shift = "0";
defparam pll7.compensate_clock = "clock0";
defparam pll7.inclk0_input_frequency = 20000;
defparam pll7.inclk1_input_frequency = 0;
defparam pll7.loop_filter_c_bits = 2;
defparam pll7.loop_filter_r_bits = 1;
defparam pll7.m = 18;
defparam pll7.m_initial = 2;
defparam pll7.m_ph = 4;
defparam pll7.n = 1;
defparam pll7.operation_mode = "normal";
defparam pll7.pfd_max = 0;
defparam pll7.pfd_min = 0;
defparam pll7.self_reset_on_loss_lock = "off";
defparam pll7.simulation_type = "timing";
defparam pll7.switch_over_type = "auto";
defparam pll7.vco_center = 0;
defparam pll7.vco_divide_by = 0;
defparam pll7.vco_frequency_control = "auto";
defparam pll7.vco_max = 0;
defparam pll7.vco_min = 0;
defparam pll7.vco_multiply_by = 0;
defparam pll7.vco_phase_shift_step = 0;
defparam pll7.vco_post_scale = 1;

cycloneive_lcell_comb locked(
	.dataa(wire_pll7_locked),
	.datab(\pll_lock_sync~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(locked1),
	.cout());
defparam locked.lut_mask = 16'hEEEE;
defparam locked.sum_lutc_input = "datac";

dffeas pll_lock_sync(
	.clk(wire_pll7_locked),
	.d(vcc),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_lock_sync~q ),
	.prn(vcc));
defparam pll_lock_sync.is_wysiwyg = "true";
defparam pll_lock_sync.power_up = "low";

endmodule

module niosII_niosII_sys_pll_stdsync_sv6 (
	altera_reset_synchronizer_int_chain_out,
	dffe6a_0,
	locked,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	dffe6a_0;
input 	locked;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosII_niosII_sys_pll_dffpipe_l2c dffpipe3(
	.clrn(altera_reset_synchronizer_int_chain_out),
	.dffe6a_0(dffe6a_0),
	.d({locked}),
	.clock(clk_clk));

endmodule

module niosII_niosII_sys_pll_dffpipe_l2c (
	clrn,
	dffe6a_0,
	d,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clrn;
output 	dffe6a_0;
input 	[0:0] d;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffe4a[0]~q ;
wire \dffe5a[0]~q ;


dffeas \dffe6a[0] (
	.clk(clock),
	.d(\dffe5a[0]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe6a_0),
	.prn(vcc));
defparam \dffe6a[0] .is_wysiwyg = "true";
defparam \dffe6a[0] .power_up = "low";

dffeas \dffe4a[0] (
	.clk(clock),
	.d(d[0]),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe4a[0]~q ),
	.prn(vcc));
defparam \dffe4a[0] .is_wysiwyg = "true";
defparam \dffe4a[0] .power_up = "low";

dffeas \dffe5a[0] (
	.clk(clock),
	.d(\dffe4a[0]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe5a[0]~q ),
	.prn(vcc));
defparam \dffe5a[0] .is_wysiwyg = "true";
defparam \dffe5a[0] .power_up = "low";

endmodule

module niosII_niosII_timer_0 (
	clk,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	reset_n,
	hold_waitrequest,
	d_write,
	write_accepted,
	read_mux_out,
	writedata,
	Equal6,
	Equal4,
	mem_used_1,
	wait_latency_counter_0,
	wait_latency_counter_1,
	Equal61,
	uav_write,
	period_l_wr_strobe1,
	timeout_occurred1,
	control_register_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_15,
	readdata_14,
	readdata_13,
	readdata_12,
	readdata_11,
	readdata_10,
	readdata_9,
	readdata_8)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	reset_n;
input 	hold_waitrequest;
input 	d_write;
input 	write_accepted;
output 	read_mux_out;
input 	[15:0] writedata;
output 	Equal6;
input 	Equal4;
input 	mem_used_1;
input 	wait_latency_counter_0;
input 	wait_latency_counter_1;
output 	Equal61;
input 	uav_write;
output 	period_l_wr_strobe1;
output 	timeout_occurred1;
output 	control_register_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_15;
output 	readdata_14;
output 	readdata_13;
output 	readdata_12;
output 	readdata_11;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \internal_counter[0]~32_combout ;
wire \period_l_register[0]~0_combout ;
wire \Equal6~2_combout ;
wire \period_l_wr_strobe~combout ;
wire \period_l_register[0]~q ;
wire \period_l_wr_strobe~3_combout ;
wire \force_reload~0_combout ;
wire \force_reload~q ;
wire \always0~0_combout ;
wire \control_wr_strobe~combout ;
wire \control_register[1]~q ;
wire \counter_is_running~0_combout ;
wire \counter_is_running~1_combout ;
wire \counter_is_running~q ;
wire \always0~1_combout ;
wire \internal_counter[0]~q ;
wire \internal_counter[0]~33 ;
wire \internal_counter[1]~34_combout ;
wire \period_l_register[1]~1_combout ;
wire \period_l_register[1]~q ;
wire \internal_counter[1]~q ;
wire \internal_counter[1]~35 ;
wire \internal_counter[2]~36_combout ;
wire \period_l_register[2]~2_combout ;
wire \period_l_register[2]~q ;
wire \internal_counter[2]~q ;
wire \internal_counter[2]~37 ;
wire \internal_counter[3]~38_combout ;
wire \period_l_register[3]~3_combout ;
wire \period_l_register[3]~q ;
wire \internal_counter[3]~q ;
wire \Equal0~0_combout ;
wire \internal_counter[3]~39 ;
wire \internal_counter[4]~40_combout ;
wire \period_l_register[4]~4_combout ;
wire \period_l_register[4]~q ;
wire \internal_counter[4]~q ;
wire \internal_counter[4]~41 ;
wire \internal_counter[5]~42_combout ;
wire \period_l_register[5]~q ;
wire \internal_counter[5]~q ;
wire \internal_counter[5]~43 ;
wire \internal_counter[6]~44_combout ;
wire \period_l_register[6]~q ;
wire \internal_counter[6]~q ;
wire \internal_counter[6]~45 ;
wire \internal_counter[7]~46_combout ;
wire \period_l_register[7]~5_combout ;
wire \period_l_register[7]~q ;
wire \internal_counter[7]~q ;
wire \Equal0~1_combout ;
wire \internal_counter[7]~47 ;
wire \internal_counter[8]~48_combout ;
wire \period_l_register[8]~q ;
wire \internal_counter[8]~q ;
wire \internal_counter[8]~49 ;
wire \internal_counter[9]~50_combout ;
wire \period_l_register[9]~6_combout ;
wire \period_l_register[9]~q ;
wire \internal_counter[9]~q ;
wire \internal_counter[9]~51 ;
wire \internal_counter[10]~52_combout ;
wire \period_l_register[10]~7_combout ;
wire \period_l_register[10]~q ;
wire \internal_counter[10]~q ;
wire \internal_counter[10]~53 ;
wire \internal_counter[11]~54_combout ;
wire \period_l_register[11]~q ;
wire \internal_counter[11]~q ;
wire \Equal0~2_combout ;
wire \internal_counter[11]~55 ;
wire \internal_counter[12]~56_combout ;
wire \period_l_register[12]~q ;
wire \internal_counter[12]~q ;
wire \internal_counter[12]~57 ;
wire \internal_counter[13]~58_combout ;
wire \period_l_register[13]~q ;
wire \internal_counter[13]~q ;
wire \internal_counter[13]~59 ;
wire \internal_counter[14]~60_combout ;
wire \period_l_register[14]~q ;
wire \internal_counter[14]~q ;
wire \internal_counter[14]~61 ;
wire \internal_counter[15]~62_combout ;
wire \period_l_register[15]~8_combout ;
wire \period_l_register[15]~q ;
wire \internal_counter[15]~q ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \internal_counter[15]~63 ;
wire \internal_counter[16]~64_combout ;
wire \period_h_register[0]~0_combout ;
wire \Equal6~3_combout ;
wire \period_h_wr_strobe~combout ;
wire \period_h_register[0]~q ;
wire \internal_counter[16]~q ;
wire \internal_counter[16]~65 ;
wire \internal_counter[17]~66_combout ;
wire \period_h_register[1]~q ;
wire \internal_counter[17]~q ;
wire \internal_counter[17]~67 ;
wire \internal_counter[18]~68_combout ;
wire \period_h_register[2]~q ;
wire \internal_counter[18]~q ;
wire \internal_counter[18]~69 ;
wire \internal_counter[19]~70_combout ;
wire \period_h_register[3]~q ;
wire \internal_counter[19]~q ;
wire \Equal0~5_combout ;
wire \internal_counter[19]~71 ;
wire \internal_counter[20]~72_combout ;
wire \period_h_register[4]~q ;
wire \internal_counter[20]~q ;
wire \internal_counter[20]~73 ;
wire \internal_counter[21]~74_combout ;
wire \period_h_register[5]~q ;
wire \internal_counter[21]~q ;
wire \internal_counter[21]~75 ;
wire \internal_counter[22]~76_combout ;
wire \period_h_register[6]~q ;
wire \internal_counter[22]~q ;
wire \internal_counter[22]~77 ;
wire \internal_counter[23]~78_combout ;
wire \period_h_register[7]~q ;
wire \internal_counter[23]~q ;
wire \Equal0~6_combout ;
wire \Equal0~7_combout ;
wire \internal_counter[23]~79 ;
wire \internal_counter[24]~80_combout ;
wire \period_h_register[8]~q ;
wire \internal_counter[24]~q ;
wire \internal_counter[24]~81 ;
wire \internal_counter[25]~82_combout ;
wire \period_h_register[9]~q ;
wire \internal_counter[25]~q ;
wire \internal_counter[25]~83 ;
wire \internal_counter[26]~84_combout ;
wire \period_h_register[10]~q ;
wire \internal_counter[26]~q ;
wire \internal_counter[26]~85 ;
wire \internal_counter[27]~86_combout ;
wire \period_h_register[11]~q ;
wire \internal_counter[27]~q ;
wire \Equal0~8_combout ;
wire \internal_counter[27]~87 ;
wire \internal_counter[28]~88_combout ;
wire \period_h_register[12]~q ;
wire \internal_counter[28]~q ;
wire \internal_counter[28]~89 ;
wire \internal_counter[29]~90_combout ;
wire \period_h_register[13]~q ;
wire \internal_counter[29]~q ;
wire \internal_counter[29]~91 ;
wire \internal_counter[30]~92_combout ;
wire \period_h_register[14]~q ;
wire \internal_counter[30]~q ;
wire \internal_counter[30]~93 ;
wire \internal_counter[31]~94_combout ;
wire \period_h_register[15]~q ;
wire \internal_counter[31]~q ;
wire \Equal0~9_combout ;
wire \Equal0~10_combout ;
wire \delayed_unxcounter_is_zeroxx0~q ;
wire \status_wr_strobe~0_combout ;
wire \timeout_occurred~0_combout ;
wire \read_mux_out[0]~1_combout ;
wire \counter_snapshot[0]~0_combout ;
wire \snap_strobe~0_combout ;
wire \counter_snapshot[0]~q ;
wire \counter_snapshot[16]~1_combout ;
wire \counter_snapshot[16]~q ;
wire \Equal6~4_combout ;
wire \Equal6~5_combout ;
wire \read_mux_out[0]~2_combout ;
wire \read_mux_out[0]~3_combout ;
wire \read_mux_out[0]~combout ;
wire \read_mux_out[1]~4_combout ;
wire \counter_snapshot[17]~q ;
wire \counter_snapshot[1]~2_combout ;
wire \counter_snapshot[1]~q ;
wire \read_mux_out[1]~5_combout ;
wire \read_mux_out[1]~6_combout ;
wire \read_mux_out[1]~combout ;
wire \read_mux_out[2]~7_combout ;
wire \counter_snapshot[18]~q ;
wire \counter_snapshot[2]~3_combout ;
wire \counter_snapshot[2]~q ;
wire \read_mux_out[2]~8_combout ;
wire \control_register[2]~q ;
wire \read_mux_out[2]~combout ;
wire \read_mux_out[3]~9_combout ;
wire \counter_snapshot[19]~q ;
wire \counter_snapshot[3]~4_combout ;
wire \counter_snapshot[3]~q ;
wire \read_mux_out[3]~10_combout ;
wire \control_register[3]~q ;
wire \read_mux_out[3]~combout ;
wire \read_mux_out[4]~11_combout ;
wire \counter_snapshot[4]~5_combout ;
wire \counter_snapshot[4]~q ;
wire \read_mux_out~12_combout ;
wire \counter_snapshot[20]~q ;
wire \read_mux_out[4]~13_combout ;
wire \read_mux_out[5]~14_combout ;
wire \counter_snapshot[5]~q ;
wire \read_mux_out~15_combout ;
wire \counter_snapshot[21]~q ;
wire \read_mux_out[5]~16_combout ;
wire \read_mux_out[6]~17_combout ;
wire \counter_snapshot[6]~q ;
wire \read_mux_out~18_combout ;
wire \counter_snapshot[22]~q ;
wire \read_mux_out[6]~19_combout ;
wire \read_mux_out[7]~20_combout ;
wire \counter_snapshot[7]~6_combout ;
wire \counter_snapshot[7]~q ;
wire \read_mux_out~21_combout ;
wire \counter_snapshot[23]~q ;
wire \read_mux_out[7]~22_combout ;
wire \read_mux_out[15]~23_combout ;
wire \counter_snapshot[15]~7_combout ;
wire \counter_snapshot[15]~q ;
wire \read_mux_out~24_combout ;
wire \counter_snapshot[31]~q ;
wire \read_mux_out[15]~25_combout ;
wire \read_mux_out[14]~26_combout ;
wire \counter_snapshot[14]~q ;
wire \read_mux_out~27_combout ;
wire \counter_snapshot[30]~q ;
wire \read_mux_out[14]~28_combout ;
wire \read_mux_out[13]~29_combout ;
wire \counter_snapshot[13]~q ;
wire \read_mux_out~30_combout ;
wire \counter_snapshot[29]~q ;
wire \read_mux_out[13]~31_combout ;
wire \read_mux_out[12]~32_combout ;
wire \counter_snapshot[12]~q ;
wire \read_mux_out~33_combout ;
wire \counter_snapshot[28]~q ;
wire \read_mux_out[12]~34_combout ;
wire \read_mux_out[11]~35_combout ;
wire \counter_snapshot[11]~q ;
wire \read_mux_out~36_combout ;
wire \counter_snapshot[27]~q ;
wire \read_mux_out[11]~37_combout ;
wire \read_mux_out[10]~38_combout ;
wire \counter_snapshot[10]~8_combout ;
wire \counter_snapshot[10]~q ;
wire \read_mux_out~39_combout ;
wire \counter_snapshot[26]~q ;
wire \read_mux_out[10]~40_combout ;
wire \read_mux_out[9]~41_combout ;
wire \counter_snapshot[9]~9_combout ;
wire \counter_snapshot[9]~q ;
wire \read_mux_out~42_combout ;
wire \counter_snapshot[25]~q ;
wire \read_mux_out[9]~43_combout ;
wire \read_mux_out[8]~44_combout ;
wire \counter_snapshot[8]~q ;
wire \read_mux_out~45_combout ;
wire \counter_snapshot[24]~q ;
wire \read_mux_out[8]~46_combout ;


cycloneive_lcell_comb \read_mux_out~0 (
	.dataa(gnd),
	.datab(W_alu_result_4),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(read_mux_out),
	.cout());
defparam \read_mux_out~0 .lut_mask = 16'h3FFF;
defparam \read_mux_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(Equal6),
	.cout());
defparam \Equal6~0 .lut_mask = 16'h0FFF;
defparam \Equal6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~1 (
	.dataa(W_alu_result_2),
	.datab(gnd),
	.datac(W_alu_result_4),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(Equal61),
	.cout());
defparam \Equal6~1 .lut_mask = 16'hAFFF;
defparam \Equal6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \period_l_wr_strobe~2 (
	.dataa(hold_waitrequest),
	.datab(Equal4),
	.datac(mem_used_1),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(period_l_wr_strobe1),
	.cout());
defparam \period_l_wr_strobe~2 .lut_mask = 16'hEFFF;
defparam \period_l_wr_strobe~2 .sum_lutc_input = "datac";

dffeas timeout_occurred(
	.clk(clk),
	.d(\timeout_occurred~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(timeout_occurred1),
	.prn(vcc));
defparam timeout_occurred.is_wysiwyg = "true";
defparam timeout_occurred.power_up = "low";

dffeas \control_register[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(control_register_0),
	.prn(vcc));
defparam \control_register[0] .is_wysiwyg = "true";
defparam \control_register[0] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk),
	.d(\read_mux_out[4]~13_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk),
	.d(\read_mux_out[5]~16_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk),
	.d(\read_mux_out[6]~19_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk),
	.d(\read_mux_out[7]~22_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk),
	.d(\read_mux_out[15]~25_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk),
	.d(\read_mux_out[14]~28_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk),
	.d(\read_mux_out[13]~31_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk),
	.d(\read_mux_out[12]~34_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk),
	.d(\read_mux_out[11]~37_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk),
	.d(\read_mux_out[10]~40_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk),
	.d(\read_mux_out[9]~43_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk),
	.d(\read_mux_out[8]~46_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

cycloneive_lcell_comb \internal_counter[0]~32 (
	.dataa(\internal_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\internal_counter[0]~32_combout ),
	.cout(\internal_counter[0]~33 ));
defparam \internal_counter[0]~32 .lut_mask = 16'h5555;
defparam \internal_counter[0]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \period_l_register[0]~0 (
	.dataa(writedata[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_l_register[0]~0_combout ),
	.cout());
defparam \period_l_register[0]~0 .lut_mask = 16'h5555;
defparam \period_l_register[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~2 (
	.dataa(W_alu_result_3),
	.datab(gnd),
	.datac(W_alu_result_4),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\Equal6~2_combout ),
	.cout());
defparam \Equal6~2 .lut_mask = 16'hAFFF;
defparam \Equal6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb period_l_wr_strobe(
	.dataa(uav_write),
	.datab(period_l_wr_strobe1),
	.datac(\Equal6~2_combout ),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\period_l_wr_strobe~combout ),
	.cout());
defparam period_l_wr_strobe.lut_mask = 16'hFEFF;
defparam period_l_wr_strobe.sum_lutc_input = "datac";

dffeas \period_l_register[0] (
	.clk(clk),
	.d(\period_l_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[0]~q ),
	.prn(vcc));
defparam \period_l_register[0] .is_wysiwyg = "true";
defparam \period_l_register[0] .power_up = "low";

cycloneive_lcell_comb \period_l_wr_strobe~3 (
	.dataa(d_write),
	.datab(write_accepted),
	.datac(period_l_wr_strobe1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\period_l_wr_strobe~3_combout ),
	.cout());
defparam \period_l_wr_strobe~3 .lut_mask = 16'hFBFF;
defparam \period_l_wr_strobe~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \force_reload~0 (
	.dataa(W_alu_result_3),
	.datab(\period_l_wr_strobe~3_combout ),
	.datac(gnd),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(\force_reload~0_combout ),
	.cout());
defparam \force_reload~0 .lut_mask = 16'hEEFF;
defparam \force_reload~0 .sum_lutc_input = "datac";

dffeas force_reload(
	.clk(clk),
	.d(\force_reload~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\force_reload~q ),
	.prn(vcc));
defparam force_reload.is_wysiwyg = "true";
defparam force_reload.power_up = "low";

cycloneive_lcell_comb \always0~0 (
	.dataa(\Equal0~10_combout ),
	.datab(\force_reload~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hEEEE;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb control_wr_strobe(
	.dataa(uav_write),
	.datab(Equal61),
	.datac(period_l_wr_strobe1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\control_wr_strobe~combout ),
	.cout());
defparam control_wr_strobe.lut_mask = 16'hFEFF;
defparam control_wr_strobe.sum_lutc_input = "datac";

dffeas \control_register[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_register[1]~q ),
	.prn(vcc));
defparam \control_register[1] .is_wysiwyg = "true";
defparam \control_register[1] .power_up = "low";

cycloneive_lcell_comb \counter_is_running~0 (
	.dataa(\counter_is_running~q ),
	.datab(\control_register[1]~q ),
	.datac(\Equal0~10_combout ),
	.datad(\force_reload~q ),
	.cin(gnd),
	.combout(\counter_is_running~0_combout ),
	.cout());
defparam \counter_is_running~0 .lut_mask = 16'hEFFF;
defparam \counter_is_running~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter_is_running~1 (
	.dataa(writedata[2]),
	.datab(\counter_is_running~0_combout ),
	.datac(\control_wr_strobe~combout ),
	.datad(writedata[3]),
	.cin(gnd),
	.combout(\counter_is_running~1_combout ),
	.cout());
defparam \counter_is_running~1 .lut_mask = 16'hACFF;
defparam \counter_is_running~1 .sum_lutc_input = "datac";

dffeas counter_is_running(
	.clk(clk),
	.d(\counter_is_running~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter_is_running~q ),
	.prn(vcc));
defparam counter_is_running.is_wysiwyg = "true";
defparam counter_is_running.power_up = "low";

cycloneive_lcell_comb \always0~1 (
	.dataa(\force_reload~q ),
	.datab(\counter_is_running~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hEEEE;
defparam \always0~1 .sum_lutc_input = "datac";

dffeas \internal_counter[0] (
	.clk(clk),
	.d(\internal_counter[0]~32_combout ),
	.asdata(\period_l_register[0]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[0]~q ),
	.prn(vcc));
defparam \internal_counter[0] .is_wysiwyg = "true";
defparam \internal_counter[0] .power_up = "low";

cycloneive_lcell_comb \internal_counter[1]~34 (
	.dataa(\internal_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[0]~33 ),
	.combout(\internal_counter[1]~34_combout ),
	.cout(\internal_counter[1]~35 ));
defparam \internal_counter[1]~34 .lut_mask = 16'h5AAF;
defparam \internal_counter[1]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \period_l_register[1]~1 (
	.dataa(writedata[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_l_register[1]~1_combout ),
	.cout());
defparam \period_l_register[1]~1 .lut_mask = 16'h5555;
defparam \period_l_register[1]~1 .sum_lutc_input = "datac";

dffeas \period_l_register[1] (
	.clk(clk),
	.d(\period_l_register[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[1]~q ),
	.prn(vcc));
defparam \period_l_register[1] .is_wysiwyg = "true";
defparam \period_l_register[1] .power_up = "low";

dffeas \internal_counter[1] (
	.clk(clk),
	.d(\internal_counter[1]~34_combout ),
	.asdata(\period_l_register[1]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[1]~q ),
	.prn(vcc));
defparam \internal_counter[1] .is_wysiwyg = "true";
defparam \internal_counter[1] .power_up = "low";

cycloneive_lcell_comb \internal_counter[2]~36 (
	.dataa(\internal_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[1]~35 ),
	.combout(\internal_counter[2]~36_combout ),
	.cout(\internal_counter[2]~37 ));
defparam \internal_counter[2]~36 .lut_mask = 16'h5A5F;
defparam \internal_counter[2]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \period_l_register[2]~2 (
	.dataa(writedata[2]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_l_register[2]~2_combout ),
	.cout());
defparam \period_l_register[2]~2 .lut_mask = 16'h5555;
defparam \period_l_register[2]~2 .sum_lutc_input = "datac";

dffeas \period_l_register[2] (
	.clk(clk),
	.d(\period_l_register[2]~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[2]~q ),
	.prn(vcc));
defparam \period_l_register[2] .is_wysiwyg = "true";
defparam \period_l_register[2] .power_up = "low";

dffeas \internal_counter[2] (
	.clk(clk),
	.d(\internal_counter[2]~36_combout ),
	.asdata(\period_l_register[2]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[2]~q ),
	.prn(vcc));
defparam \internal_counter[2] .is_wysiwyg = "true";
defparam \internal_counter[2] .power_up = "low";

cycloneive_lcell_comb \internal_counter[3]~38 (
	.dataa(\internal_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[2]~37 ),
	.combout(\internal_counter[3]~38_combout ),
	.cout(\internal_counter[3]~39 ));
defparam \internal_counter[3]~38 .lut_mask = 16'h5AAF;
defparam \internal_counter[3]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \period_l_register[3]~3 (
	.dataa(writedata[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_l_register[3]~3_combout ),
	.cout());
defparam \period_l_register[3]~3 .lut_mask = 16'h5555;
defparam \period_l_register[3]~3 .sum_lutc_input = "datac";

dffeas \period_l_register[3] (
	.clk(clk),
	.d(\period_l_register[3]~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[3]~q ),
	.prn(vcc));
defparam \period_l_register[3] .is_wysiwyg = "true";
defparam \period_l_register[3] .power_up = "low";

dffeas \internal_counter[3] (
	.clk(clk),
	.d(\internal_counter[3]~38_combout ),
	.asdata(\period_l_register[3]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[3]~q ),
	.prn(vcc));
defparam \internal_counter[3] .is_wysiwyg = "true";
defparam \internal_counter[3] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\internal_counter[0]~q ),
	.datab(\internal_counter[1]~q ),
	.datac(\internal_counter[2]~q ),
	.datad(\internal_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFFFE;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_counter[4]~40 (
	.dataa(\internal_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[3]~39 ),
	.combout(\internal_counter[4]~40_combout ),
	.cout(\internal_counter[4]~41 ));
defparam \internal_counter[4]~40 .lut_mask = 16'h5A5F;
defparam \internal_counter[4]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \period_l_register[4]~4 (
	.dataa(writedata[4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_l_register[4]~4_combout ),
	.cout());
defparam \period_l_register[4]~4 .lut_mask = 16'h5555;
defparam \period_l_register[4]~4 .sum_lutc_input = "datac";

dffeas \period_l_register[4] (
	.clk(clk),
	.d(\period_l_register[4]~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[4]~q ),
	.prn(vcc));
defparam \period_l_register[4] .is_wysiwyg = "true";
defparam \period_l_register[4] .power_up = "low";

dffeas \internal_counter[4] (
	.clk(clk),
	.d(\internal_counter[4]~40_combout ),
	.asdata(\period_l_register[4]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[4]~q ),
	.prn(vcc));
defparam \internal_counter[4] .is_wysiwyg = "true";
defparam \internal_counter[4] .power_up = "low";

cycloneive_lcell_comb \internal_counter[5]~42 (
	.dataa(\internal_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[4]~41 ),
	.combout(\internal_counter[5]~42_combout ),
	.cout(\internal_counter[5]~43 ));
defparam \internal_counter[5]~42 .lut_mask = 16'h5A5F;
defparam \internal_counter[5]~42 .sum_lutc_input = "cin";

dffeas \period_l_register[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[5]~q ),
	.prn(vcc));
defparam \period_l_register[5] .is_wysiwyg = "true";
defparam \period_l_register[5] .power_up = "low";

dffeas \internal_counter[5] (
	.clk(clk),
	.d(\internal_counter[5]~42_combout ),
	.asdata(\period_l_register[5]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[5]~q ),
	.prn(vcc));
defparam \internal_counter[5] .is_wysiwyg = "true";
defparam \internal_counter[5] .power_up = "low";

cycloneive_lcell_comb \internal_counter[6]~44 (
	.dataa(\internal_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[5]~43 ),
	.combout(\internal_counter[6]~44_combout ),
	.cout(\internal_counter[6]~45 ));
defparam \internal_counter[6]~44 .lut_mask = 16'h5AAF;
defparam \internal_counter[6]~44 .sum_lutc_input = "cin";

dffeas \period_l_register[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[6]~q ),
	.prn(vcc));
defparam \period_l_register[6] .is_wysiwyg = "true";
defparam \period_l_register[6] .power_up = "low";

dffeas \internal_counter[6] (
	.clk(clk),
	.d(\internal_counter[6]~44_combout ),
	.asdata(\period_l_register[6]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[6]~q ),
	.prn(vcc));
defparam \internal_counter[6] .is_wysiwyg = "true";
defparam \internal_counter[6] .power_up = "low";

cycloneive_lcell_comb \internal_counter[7]~46 (
	.dataa(\internal_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[6]~45 ),
	.combout(\internal_counter[7]~46_combout ),
	.cout(\internal_counter[7]~47 ));
defparam \internal_counter[7]~46 .lut_mask = 16'h5AAF;
defparam \internal_counter[7]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \period_l_register[7]~5 (
	.dataa(writedata[7]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_l_register[7]~5_combout ),
	.cout());
defparam \period_l_register[7]~5 .lut_mask = 16'h5555;
defparam \period_l_register[7]~5 .sum_lutc_input = "datac";

dffeas \period_l_register[7] (
	.clk(clk),
	.d(\period_l_register[7]~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[7]~q ),
	.prn(vcc));
defparam \period_l_register[7] .is_wysiwyg = "true";
defparam \period_l_register[7] .power_up = "low";

dffeas \internal_counter[7] (
	.clk(clk),
	.d(\internal_counter[7]~46_combout ),
	.asdata(\period_l_register[7]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[7]~q ),
	.prn(vcc));
defparam \internal_counter[7] .is_wysiwyg = "true";
defparam \internal_counter[7] .power_up = "low";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\internal_counter[4]~q ),
	.datab(\internal_counter[7]~q ),
	.datac(\internal_counter[5]~q ),
	.datad(\internal_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_counter[8]~48 (
	.dataa(\internal_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[7]~47 ),
	.combout(\internal_counter[8]~48_combout ),
	.cout(\internal_counter[8]~49 ));
defparam \internal_counter[8]~48 .lut_mask = 16'h5AAF;
defparam \internal_counter[8]~48 .sum_lutc_input = "cin";

dffeas \period_l_register[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[8]~q ),
	.prn(vcc));
defparam \period_l_register[8] .is_wysiwyg = "true";
defparam \period_l_register[8] .power_up = "low";

dffeas \internal_counter[8] (
	.clk(clk),
	.d(\internal_counter[8]~48_combout ),
	.asdata(\period_l_register[8]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[8]~q ),
	.prn(vcc));
defparam \internal_counter[8] .is_wysiwyg = "true";
defparam \internal_counter[8] .power_up = "low";

cycloneive_lcell_comb \internal_counter[9]~50 (
	.dataa(\internal_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[8]~49 ),
	.combout(\internal_counter[9]~50_combout ),
	.cout(\internal_counter[9]~51 ));
defparam \internal_counter[9]~50 .lut_mask = 16'h5AAF;
defparam \internal_counter[9]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \period_l_register[9]~6 (
	.dataa(writedata[9]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_l_register[9]~6_combout ),
	.cout());
defparam \period_l_register[9]~6 .lut_mask = 16'h5555;
defparam \period_l_register[9]~6 .sum_lutc_input = "datac";

dffeas \period_l_register[9] (
	.clk(clk),
	.d(\period_l_register[9]~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[9]~q ),
	.prn(vcc));
defparam \period_l_register[9] .is_wysiwyg = "true";
defparam \period_l_register[9] .power_up = "low";

dffeas \internal_counter[9] (
	.clk(clk),
	.d(\internal_counter[9]~50_combout ),
	.asdata(\period_l_register[9]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[9]~q ),
	.prn(vcc));
defparam \internal_counter[9] .is_wysiwyg = "true";
defparam \internal_counter[9] .power_up = "low";

cycloneive_lcell_comb \internal_counter[10]~52 (
	.dataa(\internal_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[9]~51 ),
	.combout(\internal_counter[10]~52_combout ),
	.cout(\internal_counter[10]~53 ));
defparam \internal_counter[10]~52 .lut_mask = 16'h5A5F;
defparam \internal_counter[10]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \period_l_register[10]~7 (
	.dataa(writedata[10]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_l_register[10]~7_combout ),
	.cout());
defparam \period_l_register[10]~7 .lut_mask = 16'h5555;
defparam \period_l_register[10]~7 .sum_lutc_input = "datac";

dffeas \period_l_register[10] (
	.clk(clk),
	.d(\period_l_register[10]~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[10]~q ),
	.prn(vcc));
defparam \period_l_register[10] .is_wysiwyg = "true";
defparam \period_l_register[10] .power_up = "low";

dffeas \internal_counter[10] (
	.clk(clk),
	.d(\internal_counter[10]~52_combout ),
	.asdata(\period_l_register[10]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[10]~q ),
	.prn(vcc));
defparam \internal_counter[10] .is_wysiwyg = "true";
defparam \internal_counter[10] .power_up = "low";

cycloneive_lcell_comb \internal_counter[11]~54 (
	.dataa(\internal_counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[10]~53 ),
	.combout(\internal_counter[11]~54_combout ),
	.cout(\internal_counter[11]~55 ));
defparam \internal_counter[11]~54 .lut_mask = 16'h5A5F;
defparam \internal_counter[11]~54 .sum_lutc_input = "cin";

dffeas \period_l_register[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[11]~q ),
	.prn(vcc));
defparam \period_l_register[11] .is_wysiwyg = "true";
defparam \period_l_register[11] .power_up = "low";

dffeas \internal_counter[11] (
	.clk(clk),
	.d(\internal_counter[11]~54_combout ),
	.asdata(\period_l_register[11]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[11]~q ),
	.prn(vcc));
defparam \internal_counter[11] .is_wysiwyg = "true";
defparam \internal_counter[11] .power_up = "low";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\internal_counter[9]~q ),
	.datab(\internal_counter[10]~q ),
	.datac(\internal_counter[8]~q ),
	.datad(\internal_counter[11]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEFFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_counter[12]~56 (
	.dataa(\internal_counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[11]~55 ),
	.combout(\internal_counter[12]~56_combout ),
	.cout(\internal_counter[12]~57 ));
defparam \internal_counter[12]~56 .lut_mask = 16'h5AAF;
defparam \internal_counter[12]~56 .sum_lutc_input = "cin";

dffeas \period_l_register[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[12]~q ),
	.prn(vcc));
defparam \period_l_register[12] .is_wysiwyg = "true";
defparam \period_l_register[12] .power_up = "low";

dffeas \internal_counter[12] (
	.clk(clk),
	.d(\internal_counter[12]~56_combout ),
	.asdata(\period_l_register[12]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[12]~q ),
	.prn(vcc));
defparam \internal_counter[12] .is_wysiwyg = "true";
defparam \internal_counter[12] .power_up = "low";

cycloneive_lcell_comb \internal_counter[13]~58 (
	.dataa(\internal_counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[12]~57 ),
	.combout(\internal_counter[13]~58_combout ),
	.cout(\internal_counter[13]~59 ));
defparam \internal_counter[13]~58 .lut_mask = 16'h5A5F;
defparam \internal_counter[13]~58 .sum_lutc_input = "cin";

dffeas \period_l_register[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[13]~q ),
	.prn(vcc));
defparam \period_l_register[13] .is_wysiwyg = "true";
defparam \period_l_register[13] .power_up = "low";

dffeas \internal_counter[13] (
	.clk(clk),
	.d(\internal_counter[13]~58_combout ),
	.asdata(\period_l_register[13]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[13]~q ),
	.prn(vcc));
defparam \internal_counter[13] .is_wysiwyg = "true";
defparam \internal_counter[13] .power_up = "low";

cycloneive_lcell_comb \internal_counter[14]~60 (
	.dataa(\internal_counter[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[13]~59 ),
	.combout(\internal_counter[14]~60_combout ),
	.cout(\internal_counter[14]~61 ));
defparam \internal_counter[14]~60 .lut_mask = 16'h5AAF;
defparam \internal_counter[14]~60 .sum_lutc_input = "cin";

dffeas \period_l_register[14] (
	.clk(clk),
	.d(writedata[14]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[14]~q ),
	.prn(vcc));
defparam \period_l_register[14] .is_wysiwyg = "true";
defparam \period_l_register[14] .power_up = "low";

dffeas \internal_counter[14] (
	.clk(clk),
	.d(\internal_counter[14]~60_combout ),
	.asdata(\period_l_register[14]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[14]~q ),
	.prn(vcc));
defparam \internal_counter[14] .is_wysiwyg = "true";
defparam \internal_counter[14] .power_up = "low";

cycloneive_lcell_comb \internal_counter[15]~62 (
	.dataa(\internal_counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[14]~61 ),
	.combout(\internal_counter[15]~62_combout ),
	.cout(\internal_counter[15]~63 ));
defparam \internal_counter[15]~62 .lut_mask = 16'h5AAF;
defparam \internal_counter[15]~62 .sum_lutc_input = "cin";

cycloneive_lcell_comb \period_l_register[15]~8 (
	.dataa(writedata[15]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_l_register[15]~8_combout ),
	.cout());
defparam \period_l_register[15]~8 .lut_mask = 16'h5555;
defparam \period_l_register[15]~8 .sum_lutc_input = "datac";

dffeas \period_l_register[15] (
	.clk(clk),
	.d(\period_l_register[15]~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[15]~q ),
	.prn(vcc));
defparam \period_l_register[15] .is_wysiwyg = "true";
defparam \period_l_register[15] .power_up = "low";

dffeas \internal_counter[15] (
	.clk(clk),
	.d(\internal_counter[15]~62_combout ),
	.asdata(\period_l_register[15]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[15]~q ),
	.prn(vcc));
defparam \internal_counter[15] .is_wysiwyg = "true";
defparam \internal_counter[15] .power_up = "low";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\internal_counter[15]~q ),
	.datab(\internal_counter[12]~q ),
	.datac(\internal_counter[13]~q ),
	.datad(\internal_counter[14]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hBFFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'hFFFE;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_counter[16]~64 (
	.dataa(\internal_counter[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[15]~63 ),
	.combout(\internal_counter[16]~64_combout ),
	.cout(\internal_counter[16]~65 ));
defparam \internal_counter[16]~64 .lut_mask = 16'h5A5F;
defparam \internal_counter[16]~64 .sum_lutc_input = "cin";

cycloneive_lcell_comb \period_h_register[0]~0 (
	.dataa(writedata[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\period_h_register[0]~0_combout ),
	.cout());
defparam \period_h_register[0]~0 .lut_mask = 16'h5555;
defparam \period_h_register[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~3 (
	.dataa(W_alu_result_3),
	.datab(W_alu_result_2),
	.datac(gnd),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(\Equal6~3_combout ),
	.cout());
defparam \Equal6~3 .lut_mask = 16'hEEFF;
defparam \Equal6~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb period_h_wr_strobe(
	.dataa(uav_write),
	.datab(period_l_wr_strobe1),
	.datac(\Equal6~3_combout ),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\period_h_wr_strobe~combout ),
	.cout());
defparam period_h_wr_strobe.lut_mask = 16'hFEFF;
defparam period_h_wr_strobe.sum_lutc_input = "datac";

dffeas \period_h_register[0] (
	.clk(clk),
	.d(\period_h_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[0]~q ),
	.prn(vcc));
defparam \period_h_register[0] .is_wysiwyg = "true";
defparam \period_h_register[0] .power_up = "low";

dffeas \internal_counter[16] (
	.clk(clk),
	.d(\internal_counter[16]~64_combout ),
	.asdata(\period_h_register[0]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[16]~q ),
	.prn(vcc));
defparam \internal_counter[16] .is_wysiwyg = "true";
defparam \internal_counter[16] .power_up = "low";

cycloneive_lcell_comb \internal_counter[17]~66 (
	.dataa(\internal_counter[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[16]~65 ),
	.combout(\internal_counter[17]~66_combout ),
	.cout(\internal_counter[17]~67 ));
defparam \internal_counter[17]~66 .lut_mask = 16'h5A5F;
defparam \internal_counter[17]~66 .sum_lutc_input = "cin";

dffeas \period_h_register[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[1]~q ),
	.prn(vcc));
defparam \period_h_register[1] .is_wysiwyg = "true";
defparam \period_h_register[1] .power_up = "low";

dffeas \internal_counter[17] (
	.clk(clk),
	.d(\internal_counter[17]~66_combout ),
	.asdata(\period_h_register[1]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[17]~q ),
	.prn(vcc));
defparam \internal_counter[17] .is_wysiwyg = "true";
defparam \internal_counter[17] .power_up = "low";

cycloneive_lcell_comb \internal_counter[18]~68 (
	.dataa(\internal_counter[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[17]~67 ),
	.combout(\internal_counter[18]~68_combout ),
	.cout(\internal_counter[18]~69 ));
defparam \internal_counter[18]~68 .lut_mask = 16'h5AAF;
defparam \internal_counter[18]~68 .sum_lutc_input = "cin";

dffeas \period_h_register[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[2]~q ),
	.prn(vcc));
defparam \period_h_register[2] .is_wysiwyg = "true";
defparam \period_h_register[2] .power_up = "low";

dffeas \internal_counter[18] (
	.clk(clk),
	.d(\internal_counter[18]~68_combout ),
	.asdata(\period_h_register[2]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[18]~q ),
	.prn(vcc));
defparam \internal_counter[18] .is_wysiwyg = "true";
defparam \internal_counter[18] .power_up = "low";

cycloneive_lcell_comb \internal_counter[19]~70 (
	.dataa(\internal_counter[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[18]~69 ),
	.combout(\internal_counter[19]~70_combout ),
	.cout(\internal_counter[19]~71 ));
defparam \internal_counter[19]~70 .lut_mask = 16'h5A5F;
defparam \internal_counter[19]~70 .sum_lutc_input = "cin";

dffeas \period_h_register[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[3]~q ),
	.prn(vcc));
defparam \period_h_register[3] .is_wysiwyg = "true";
defparam \period_h_register[3] .power_up = "low";

dffeas \internal_counter[19] (
	.clk(clk),
	.d(\internal_counter[19]~70_combout ),
	.asdata(\period_h_register[3]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[19]~q ),
	.prn(vcc));
defparam \internal_counter[19] .is_wysiwyg = "true";
defparam \internal_counter[19] .power_up = "low";

cycloneive_lcell_comb \Equal0~5 (
	.dataa(\internal_counter[16]~q ),
	.datab(\internal_counter[17]~q ),
	.datac(\internal_counter[18]~q ),
	.datad(\internal_counter[19]~q ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'hBFFF;
defparam \Equal0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_counter[20]~72 (
	.dataa(\internal_counter[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[19]~71 ),
	.combout(\internal_counter[20]~72_combout ),
	.cout(\internal_counter[20]~73 ));
defparam \internal_counter[20]~72 .lut_mask = 16'h5AAF;
defparam \internal_counter[20]~72 .sum_lutc_input = "cin";

dffeas \period_h_register[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[4]~q ),
	.prn(vcc));
defparam \period_h_register[4] .is_wysiwyg = "true";
defparam \period_h_register[4] .power_up = "low";

dffeas \internal_counter[20] (
	.clk(clk),
	.d(\internal_counter[20]~72_combout ),
	.asdata(\period_h_register[4]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[20]~q ),
	.prn(vcc));
defparam \internal_counter[20] .is_wysiwyg = "true";
defparam \internal_counter[20] .power_up = "low";

cycloneive_lcell_comb \internal_counter[21]~74 (
	.dataa(\internal_counter[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[20]~73 ),
	.combout(\internal_counter[21]~74_combout ),
	.cout(\internal_counter[21]~75 ));
defparam \internal_counter[21]~74 .lut_mask = 16'h5A5F;
defparam \internal_counter[21]~74 .sum_lutc_input = "cin";

dffeas \period_h_register[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[5]~q ),
	.prn(vcc));
defparam \period_h_register[5] .is_wysiwyg = "true";
defparam \period_h_register[5] .power_up = "low";

dffeas \internal_counter[21] (
	.clk(clk),
	.d(\internal_counter[21]~74_combout ),
	.asdata(\period_h_register[5]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[21]~q ),
	.prn(vcc));
defparam \internal_counter[21] .is_wysiwyg = "true";
defparam \internal_counter[21] .power_up = "low";

cycloneive_lcell_comb \internal_counter[22]~76 (
	.dataa(\internal_counter[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[21]~75 ),
	.combout(\internal_counter[22]~76_combout ),
	.cout(\internal_counter[22]~77 ));
defparam \internal_counter[22]~76 .lut_mask = 16'h5AAF;
defparam \internal_counter[22]~76 .sum_lutc_input = "cin";

dffeas \period_h_register[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[6]~q ),
	.prn(vcc));
defparam \period_h_register[6] .is_wysiwyg = "true";
defparam \period_h_register[6] .power_up = "low";

dffeas \internal_counter[22] (
	.clk(clk),
	.d(\internal_counter[22]~76_combout ),
	.asdata(\period_h_register[6]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[22]~q ),
	.prn(vcc));
defparam \internal_counter[22] .is_wysiwyg = "true";
defparam \internal_counter[22] .power_up = "low";

cycloneive_lcell_comb \internal_counter[23]~78 (
	.dataa(\internal_counter[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[22]~77 ),
	.combout(\internal_counter[23]~78_combout ),
	.cout(\internal_counter[23]~79 ));
defparam \internal_counter[23]~78 .lut_mask = 16'h5A5F;
defparam \internal_counter[23]~78 .sum_lutc_input = "cin";

dffeas \period_h_register[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[7]~q ),
	.prn(vcc));
defparam \period_h_register[7] .is_wysiwyg = "true";
defparam \period_h_register[7] .power_up = "low";

dffeas \internal_counter[23] (
	.clk(clk),
	.d(\internal_counter[23]~78_combout ),
	.asdata(\period_h_register[7]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[23]~q ),
	.prn(vcc));
defparam \internal_counter[23] .is_wysiwyg = "true";
defparam \internal_counter[23] .power_up = "low";

cycloneive_lcell_comb \Equal0~6 (
	.dataa(\internal_counter[20]~q ),
	.datab(\internal_counter[21]~q ),
	.datac(\internal_counter[22]~q ),
	.datad(\internal_counter[23]~q ),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
defparam \Equal0~6 .lut_mask = 16'h7FFF;
defparam \Equal0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~7 (
	.dataa(\Equal0~5_combout ),
	.datab(\Equal0~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
defparam \Equal0~7 .lut_mask = 16'hEEEE;
defparam \Equal0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_counter[24]~80 (
	.dataa(\internal_counter[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[23]~79 ),
	.combout(\internal_counter[24]~80_combout ),
	.cout(\internal_counter[24]~81 ));
defparam \internal_counter[24]~80 .lut_mask = 16'h5AAF;
defparam \internal_counter[24]~80 .sum_lutc_input = "cin";

dffeas \period_h_register[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[8]~q ),
	.prn(vcc));
defparam \period_h_register[8] .is_wysiwyg = "true";
defparam \period_h_register[8] .power_up = "low";

dffeas \internal_counter[24] (
	.clk(clk),
	.d(\internal_counter[24]~80_combout ),
	.asdata(\period_h_register[8]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[24]~q ),
	.prn(vcc));
defparam \internal_counter[24] .is_wysiwyg = "true";
defparam \internal_counter[24] .power_up = "low";

cycloneive_lcell_comb \internal_counter[25]~82 (
	.dataa(\internal_counter[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[24]~81 ),
	.combout(\internal_counter[25]~82_combout ),
	.cout(\internal_counter[25]~83 ));
defparam \internal_counter[25]~82 .lut_mask = 16'h5A5F;
defparam \internal_counter[25]~82 .sum_lutc_input = "cin";

dffeas \period_h_register[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[9]~q ),
	.prn(vcc));
defparam \period_h_register[9] .is_wysiwyg = "true";
defparam \period_h_register[9] .power_up = "low";

dffeas \internal_counter[25] (
	.clk(clk),
	.d(\internal_counter[25]~82_combout ),
	.asdata(\period_h_register[9]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[25]~q ),
	.prn(vcc));
defparam \internal_counter[25] .is_wysiwyg = "true";
defparam \internal_counter[25] .power_up = "low";

cycloneive_lcell_comb \internal_counter[26]~84 (
	.dataa(\internal_counter[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[25]~83 ),
	.combout(\internal_counter[26]~84_combout ),
	.cout(\internal_counter[26]~85 ));
defparam \internal_counter[26]~84 .lut_mask = 16'h5AAF;
defparam \internal_counter[26]~84 .sum_lutc_input = "cin";

dffeas \period_h_register[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[10]~q ),
	.prn(vcc));
defparam \period_h_register[10] .is_wysiwyg = "true";
defparam \period_h_register[10] .power_up = "low";

dffeas \internal_counter[26] (
	.clk(clk),
	.d(\internal_counter[26]~84_combout ),
	.asdata(\period_h_register[10]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[26]~q ),
	.prn(vcc));
defparam \internal_counter[26] .is_wysiwyg = "true";
defparam \internal_counter[26] .power_up = "low";

cycloneive_lcell_comb \internal_counter[27]~86 (
	.dataa(\internal_counter[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[26]~85 ),
	.combout(\internal_counter[27]~86_combout ),
	.cout(\internal_counter[27]~87 ));
defparam \internal_counter[27]~86 .lut_mask = 16'h5A5F;
defparam \internal_counter[27]~86 .sum_lutc_input = "cin";

dffeas \period_h_register[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[11]~q ),
	.prn(vcc));
defparam \period_h_register[11] .is_wysiwyg = "true";
defparam \period_h_register[11] .power_up = "low";

dffeas \internal_counter[27] (
	.clk(clk),
	.d(\internal_counter[27]~86_combout ),
	.asdata(\period_h_register[11]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[27]~q ),
	.prn(vcc));
defparam \internal_counter[27] .is_wysiwyg = "true";
defparam \internal_counter[27] .power_up = "low";

cycloneive_lcell_comb \Equal0~8 (
	.dataa(\internal_counter[24]~q ),
	.datab(\internal_counter[25]~q ),
	.datac(\internal_counter[26]~q ),
	.datad(\internal_counter[27]~q ),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
defparam \Equal0~8 .lut_mask = 16'h7FFF;
defparam \Equal0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_counter[28]~88 (
	.dataa(\internal_counter[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[27]~87 ),
	.combout(\internal_counter[28]~88_combout ),
	.cout(\internal_counter[28]~89 ));
defparam \internal_counter[28]~88 .lut_mask = 16'h5AAF;
defparam \internal_counter[28]~88 .sum_lutc_input = "cin";

dffeas \period_h_register[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[12]~q ),
	.prn(vcc));
defparam \period_h_register[12] .is_wysiwyg = "true";
defparam \period_h_register[12] .power_up = "low";

dffeas \internal_counter[28] (
	.clk(clk),
	.d(\internal_counter[28]~88_combout ),
	.asdata(\period_h_register[12]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[28]~q ),
	.prn(vcc));
defparam \internal_counter[28] .is_wysiwyg = "true";
defparam \internal_counter[28] .power_up = "low";

cycloneive_lcell_comb \internal_counter[29]~90 (
	.dataa(\internal_counter[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[28]~89 ),
	.combout(\internal_counter[29]~90_combout ),
	.cout(\internal_counter[29]~91 ));
defparam \internal_counter[29]~90 .lut_mask = 16'h5A5F;
defparam \internal_counter[29]~90 .sum_lutc_input = "cin";

dffeas \period_h_register[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[13]~q ),
	.prn(vcc));
defparam \period_h_register[13] .is_wysiwyg = "true";
defparam \period_h_register[13] .power_up = "low";

dffeas \internal_counter[29] (
	.clk(clk),
	.d(\internal_counter[29]~90_combout ),
	.asdata(\period_h_register[13]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[29]~q ),
	.prn(vcc));
defparam \internal_counter[29] .is_wysiwyg = "true";
defparam \internal_counter[29] .power_up = "low";

cycloneive_lcell_comb \internal_counter[30]~92 (
	.dataa(\internal_counter[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\internal_counter[29]~91 ),
	.combout(\internal_counter[30]~92_combout ),
	.cout(\internal_counter[30]~93 ));
defparam \internal_counter[30]~92 .lut_mask = 16'h5AAF;
defparam \internal_counter[30]~92 .sum_lutc_input = "cin";

dffeas \period_h_register[14] (
	.clk(clk),
	.d(writedata[14]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[14]~q ),
	.prn(vcc));
defparam \period_h_register[14] .is_wysiwyg = "true";
defparam \period_h_register[14] .power_up = "low";

dffeas \internal_counter[30] (
	.clk(clk),
	.d(\internal_counter[30]~92_combout ),
	.asdata(\period_h_register[14]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[30]~q ),
	.prn(vcc));
defparam \internal_counter[30] .is_wysiwyg = "true";
defparam \internal_counter[30] .power_up = "low";

cycloneive_lcell_comb \internal_counter[31]~94 (
	.dataa(\internal_counter[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\internal_counter[30]~93 ),
	.combout(\internal_counter[31]~94_combout ),
	.cout());
defparam \internal_counter[31]~94 .lut_mask = 16'h5A5A;
defparam \internal_counter[31]~94 .sum_lutc_input = "cin";

dffeas \period_h_register[15] (
	.clk(clk),
	.d(writedata[15]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[15]~q ),
	.prn(vcc));
defparam \period_h_register[15] .is_wysiwyg = "true";
defparam \period_h_register[15] .power_up = "low";

dffeas \internal_counter[31] (
	.clk(clk),
	.d(\internal_counter[31]~94_combout ),
	.asdata(\period_h_register[15]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[31]~q ),
	.prn(vcc));
defparam \internal_counter[31] .is_wysiwyg = "true";
defparam \internal_counter[31] .power_up = "low";

cycloneive_lcell_comb \Equal0~9 (
	.dataa(\internal_counter[28]~q ),
	.datab(\internal_counter[29]~q ),
	.datac(\internal_counter[30]~q ),
	.datad(\internal_counter[31]~q ),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
defparam \Equal0~9 .lut_mask = 16'h7FFF;
defparam \Equal0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~10 (
	.dataa(\Equal0~4_combout ),
	.datab(\Equal0~7_combout ),
	.datac(\Equal0~8_combout ),
	.datad(\Equal0~9_combout ),
	.cin(gnd),
	.combout(\Equal0~10_combout ),
	.cout());
defparam \Equal0~10 .lut_mask = 16'hFFFE;
defparam \Equal0~10 .sum_lutc_input = "datac";

dffeas delayed_unxcounter_is_zeroxx0(
	.clk(clk),
	.d(\Equal0~10_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_unxcounter_is_zeroxx0~q ),
	.prn(vcc));
defparam delayed_unxcounter_is_zeroxx0.is_wysiwyg = "true";
defparam delayed_unxcounter_is_zeroxx0.power_up = "low";

cycloneive_lcell_comb \status_wr_strobe~0 (
	.dataa(uav_write),
	.datab(read_mux_out),
	.datac(period_l_wr_strobe1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\status_wr_strobe~0_combout ),
	.cout());
defparam \status_wr_strobe~0 .lut_mask = 16'hFEFF;
defparam \status_wr_strobe~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \timeout_occurred~0 (
	.dataa(timeout_occurred1),
	.datab(\Equal0~10_combout ),
	.datac(\delayed_unxcounter_is_zeroxx0~q ),
	.datad(\status_wr_strobe~0_combout ),
	.cin(gnd),
	.combout(\timeout_occurred~0_combout ),
	.cout());
defparam \timeout_occurred~0 .lut_mask = 16'hEFFF;
defparam \timeout_occurred~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[0]~1 (
	.dataa(\Equal6~2_combout ),
	.datab(\Equal6~3_combout ),
	.datac(\period_l_register[0]~q ),
	.datad(\period_h_register[0]~q ),
	.cin(gnd),
	.combout(\read_mux_out[0]~1_combout ),
	.cout());
defparam \read_mux_out[0]~1 .lut_mask = 16'hEFFF;
defparam \read_mux_out[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter_snapshot[0]~0 (
	.dataa(\internal_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[0]~0_combout ),
	.cout());
defparam \counter_snapshot[0]~0 .lut_mask = 16'h5555;
defparam \counter_snapshot[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \snap_strobe~0 (
	.dataa(W_alu_result_4),
	.datab(\period_l_wr_strobe~3_combout ),
	.datac(gnd),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\snap_strobe~0_combout ),
	.cout());
defparam \snap_strobe~0 .lut_mask = 16'hEEFF;
defparam \snap_strobe~0 .sum_lutc_input = "datac";

dffeas \counter_snapshot[0] (
	.clk(clk),
	.d(\counter_snapshot[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[0]~q ),
	.prn(vcc));
defparam \counter_snapshot[0] .is_wysiwyg = "true";
defparam \counter_snapshot[0] .power_up = "low";

cycloneive_lcell_comb \counter_snapshot[16]~1 (
	.dataa(\internal_counter[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[16]~1_combout ),
	.cout());
defparam \counter_snapshot[16]~1 .lut_mask = 16'h5555;
defparam \counter_snapshot[16]~1 .sum_lutc_input = "datac";

dffeas \counter_snapshot[16] (
	.clk(clk),
	.d(\counter_snapshot[16]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[16]~q ),
	.prn(vcc));
defparam \counter_snapshot[16] .is_wysiwyg = "true";
defparam \counter_snapshot[16] .power_up = "low";

cycloneive_lcell_comb \Equal6~4 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_2),
	.datac(gnd),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\Equal6~4_combout ),
	.cout());
defparam \Equal6~4 .lut_mask = 16'hEEFF;
defparam \Equal6~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~5 (
	.dataa(W_alu_result_4),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\Equal6~5_combout ),
	.cout());
defparam \Equal6~5 .lut_mask = 16'hAFFF;
defparam \Equal6~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[0]~2 (
	.dataa(\counter_snapshot[0]~q ),
	.datab(\counter_snapshot[16]~q ),
	.datac(\Equal6~4_combout ),
	.datad(\Equal6~5_combout ),
	.cin(gnd),
	.combout(\read_mux_out[0]~2_combout ),
	.cout());
defparam \read_mux_out[0]~2 .lut_mask = 16'hFFFE;
defparam \read_mux_out[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[0]~3 (
	.dataa(read_mux_out),
	.datab(Equal61),
	.datac(control_register_0),
	.datad(timeout_occurred1),
	.cin(gnd),
	.combout(\read_mux_out[0]~3_combout ),
	.cout());
defparam \read_mux_out[0]~3 .lut_mask = 16'hFFFE;
defparam \read_mux_out[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[0] (
	.dataa(\read_mux_out[0]~1_combout ),
	.datab(\read_mux_out[0]~2_combout ),
	.datac(\read_mux_out[0]~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_mux_out[0]~combout ),
	.cout());
defparam \read_mux_out[0] .lut_mask = 16'hFEFE;
defparam \read_mux_out[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[1]~4 (
	.dataa(\Equal6~3_combout ),
	.datab(\period_h_register[1]~q ),
	.datac(\Equal6~2_combout ),
	.datad(\period_l_register[1]~q ),
	.cin(gnd),
	.combout(\read_mux_out[1]~4_combout ),
	.cout());
defparam \read_mux_out[1]~4 .lut_mask = 16'hFEFF;
defparam \read_mux_out[1]~4 .sum_lutc_input = "datac";

dffeas \counter_snapshot[17] (
	.clk(clk),
	.d(\internal_counter[17]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[17]~q ),
	.prn(vcc));
defparam \counter_snapshot[17] .is_wysiwyg = "true";
defparam \counter_snapshot[17] .power_up = "low";

cycloneive_lcell_comb \counter_snapshot[1]~2 (
	.dataa(\internal_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[1]~2_combout ),
	.cout());
defparam \counter_snapshot[1]~2 .lut_mask = 16'h5555;
defparam \counter_snapshot[1]~2 .sum_lutc_input = "datac";

dffeas \counter_snapshot[1] (
	.clk(clk),
	.d(\counter_snapshot[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[1]~q ),
	.prn(vcc));
defparam \counter_snapshot[1] .is_wysiwyg = "true";
defparam \counter_snapshot[1] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[1]~5 (
	.dataa(\Equal6~5_combout ),
	.datab(\Equal6~4_combout ),
	.datac(\counter_snapshot[17]~q ),
	.datad(\counter_snapshot[1]~q ),
	.cin(gnd),
	.combout(\read_mux_out[1]~5_combout ),
	.cout());
defparam \read_mux_out[1]~5 .lut_mask = 16'hFFFE;
defparam \read_mux_out[1]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[1]~6 (
	.dataa(read_mux_out),
	.datab(Equal61),
	.datac(\control_register[1]~q ),
	.datad(\counter_is_running~q ),
	.cin(gnd),
	.combout(\read_mux_out[1]~6_combout ),
	.cout());
defparam \read_mux_out[1]~6 .lut_mask = 16'hFFFE;
defparam \read_mux_out[1]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[1] (
	.dataa(\read_mux_out[1]~4_combout ),
	.datab(\read_mux_out[1]~5_combout ),
	.datac(\read_mux_out[1]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_mux_out[1]~combout ),
	.cout());
defparam \read_mux_out[1] .lut_mask = 16'hFEFE;
defparam \read_mux_out[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[2]~7 (
	.dataa(\Equal6~3_combout ),
	.datab(\period_h_register[2]~q ),
	.datac(\Equal6~2_combout ),
	.datad(\period_l_register[2]~q ),
	.cin(gnd),
	.combout(\read_mux_out[2]~7_combout ),
	.cout());
defparam \read_mux_out[2]~7 .lut_mask = 16'hFEFF;
defparam \read_mux_out[2]~7 .sum_lutc_input = "datac";

dffeas \counter_snapshot[18] (
	.clk(clk),
	.d(\internal_counter[18]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[18]~q ),
	.prn(vcc));
defparam \counter_snapshot[18] .is_wysiwyg = "true";
defparam \counter_snapshot[18] .power_up = "low";

cycloneive_lcell_comb \counter_snapshot[2]~3 (
	.dataa(\internal_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[2]~3_combout ),
	.cout());
defparam \counter_snapshot[2]~3 .lut_mask = 16'h5555;
defparam \counter_snapshot[2]~3 .sum_lutc_input = "datac";

dffeas \counter_snapshot[2] (
	.clk(clk),
	.d(\counter_snapshot[2]~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[2]~q ),
	.prn(vcc));
defparam \counter_snapshot[2] .is_wysiwyg = "true";
defparam \counter_snapshot[2] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[2]~8 (
	.dataa(\Equal6~5_combout ),
	.datab(\Equal6~4_combout ),
	.datac(\counter_snapshot[18]~q ),
	.datad(\counter_snapshot[2]~q ),
	.cin(gnd),
	.combout(\read_mux_out[2]~8_combout ),
	.cout());
defparam \read_mux_out[2]~8 .lut_mask = 16'hFFFE;
defparam \read_mux_out[2]~8 .sum_lutc_input = "datac";

dffeas \control_register[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_register[2]~q ),
	.prn(vcc));
defparam \control_register[2] .is_wysiwyg = "true";
defparam \control_register[2] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[2] (
	.dataa(\read_mux_out[2]~7_combout ),
	.datab(\read_mux_out[2]~8_combout ),
	.datac(Equal61),
	.datad(\control_register[2]~q ),
	.cin(gnd),
	.combout(\read_mux_out[2]~combout ),
	.cout());
defparam \read_mux_out[2] .lut_mask = 16'hFFFE;
defparam \read_mux_out[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[3]~9 (
	.dataa(\Equal6~3_combout ),
	.datab(\period_h_register[3]~q ),
	.datac(\Equal6~2_combout ),
	.datad(\period_l_register[3]~q ),
	.cin(gnd),
	.combout(\read_mux_out[3]~9_combout ),
	.cout());
defparam \read_mux_out[3]~9 .lut_mask = 16'hFEFF;
defparam \read_mux_out[3]~9 .sum_lutc_input = "datac";

dffeas \counter_snapshot[19] (
	.clk(clk),
	.d(\internal_counter[19]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[19]~q ),
	.prn(vcc));
defparam \counter_snapshot[19] .is_wysiwyg = "true";
defparam \counter_snapshot[19] .power_up = "low";

cycloneive_lcell_comb \counter_snapshot[3]~4 (
	.dataa(\internal_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[3]~4_combout ),
	.cout());
defparam \counter_snapshot[3]~4 .lut_mask = 16'h5555;
defparam \counter_snapshot[3]~4 .sum_lutc_input = "datac";

dffeas \counter_snapshot[3] (
	.clk(clk),
	.d(\counter_snapshot[3]~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[3]~q ),
	.prn(vcc));
defparam \counter_snapshot[3] .is_wysiwyg = "true";
defparam \counter_snapshot[3] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[3]~10 (
	.dataa(\Equal6~5_combout ),
	.datab(\Equal6~4_combout ),
	.datac(\counter_snapshot[19]~q ),
	.datad(\counter_snapshot[3]~q ),
	.cin(gnd),
	.combout(\read_mux_out[3]~10_combout ),
	.cout());
defparam \read_mux_out[3]~10 .lut_mask = 16'hFFFE;
defparam \read_mux_out[3]~10 .sum_lutc_input = "datac";

dffeas \control_register[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_register[3]~q ),
	.prn(vcc));
defparam \control_register[3] .is_wysiwyg = "true";
defparam \control_register[3] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[3] (
	.dataa(\read_mux_out[3]~9_combout ),
	.datab(\read_mux_out[3]~10_combout ),
	.datac(Equal61),
	.datad(\control_register[3]~q ),
	.cin(gnd),
	.combout(\read_mux_out[3]~combout ),
	.cout());
defparam \read_mux_out[3] .lut_mask = 16'hFFFE;
defparam \read_mux_out[3] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[4]~11 (
	.dataa(\Equal6~3_combout ),
	.datab(\period_h_register[4]~q ),
	.datac(\Equal6~2_combout ),
	.datad(\period_l_register[4]~q ),
	.cin(gnd),
	.combout(\read_mux_out[4]~11_combout ),
	.cout());
defparam \read_mux_out[4]~11 .lut_mask = 16'hFEFF;
defparam \read_mux_out[4]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter_snapshot[4]~5 (
	.dataa(\internal_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[4]~5_combout ),
	.cout());
defparam \counter_snapshot[4]~5 .lut_mask = 16'h5555;
defparam \counter_snapshot[4]~5 .sum_lutc_input = "datac";

dffeas \counter_snapshot[4] (
	.clk(clk),
	.d(\counter_snapshot[4]~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[4]~q ),
	.prn(vcc));
defparam \counter_snapshot[4] .is_wysiwyg = "true";
defparam \counter_snapshot[4] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~12 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[4]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~12_combout ),
	.cout());
defparam \read_mux_out~12 .lut_mask = 16'hEFFF;
defparam \read_mux_out~12 .sum_lutc_input = "datac";

dffeas \counter_snapshot[20] (
	.clk(clk),
	.d(\internal_counter[20]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[20]~q ),
	.prn(vcc));
defparam \counter_snapshot[20] .is_wysiwyg = "true";
defparam \counter_snapshot[20] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[4]~13 (
	.dataa(\read_mux_out[4]~11_combout ),
	.datab(\read_mux_out~12_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[20]~q ),
	.cin(gnd),
	.combout(\read_mux_out[4]~13_combout ),
	.cout());
defparam \read_mux_out[4]~13 .lut_mask = 16'hFFFE;
defparam \read_mux_out[4]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[5]~14 (
	.dataa(\Equal6~2_combout ),
	.datab(\Equal6~3_combout ),
	.datac(\period_h_register[5]~q ),
	.datad(\period_l_register[5]~q ),
	.cin(gnd),
	.combout(\read_mux_out[5]~14_combout ),
	.cout());
defparam \read_mux_out[5]~14 .lut_mask = 16'hFFFE;
defparam \read_mux_out[5]~14 .sum_lutc_input = "datac";

dffeas \counter_snapshot[5] (
	.clk(clk),
	.d(\internal_counter[5]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[5]~q ),
	.prn(vcc));
defparam \counter_snapshot[5] .is_wysiwyg = "true";
defparam \counter_snapshot[5] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~15 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[5]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~15_combout ),
	.cout());
defparam \read_mux_out~15 .lut_mask = 16'hEFFF;
defparam \read_mux_out~15 .sum_lutc_input = "datac";

dffeas \counter_snapshot[21] (
	.clk(clk),
	.d(\internal_counter[21]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[21]~q ),
	.prn(vcc));
defparam \counter_snapshot[21] .is_wysiwyg = "true";
defparam \counter_snapshot[21] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[5]~16 (
	.dataa(\read_mux_out[5]~14_combout ),
	.datab(\read_mux_out~15_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[21]~q ),
	.cin(gnd),
	.combout(\read_mux_out[5]~16_combout ),
	.cout());
defparam \read_mux_out[5]~16 .lut_mask = 16'hFFFE;
defparam \read_mux_out[5]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[6]~17 (
	.dataa(\Equal6~2_combout ),
	.datab(\Equal6~3_combout ),
	.datac(\period_h_register[6]~q ),
	.datad(\period_l_register[6]~q ),
	.cin(gnd),
	.combout(\read_mux_out[6]~17_combout ),
	.cout());
defparam \read_mux_out[6]~17 .lut_mask = 16'hFFFE;
defparam \read_mux_out[6]~17 .sum_lutc_input = "datac";

dffeas \counter_snapshot[6] (
	.clk(clk),
	.d(\internal_counter[6]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[6]~q ),
	.prn(vcc));
defparam \counter_snapshot[6] .is_wysiwyg = "true";
defparam \counter_snapshot[6] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~18 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[6]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~18_combout ),
	.cout());
defparam \read_mux_out~18 .lut_mask = 16'hEFFF;
defparam \read_mux_out~18 .sum_lutc_input = "datac";

dffeas \counter_snapshot[22] (
	.clk(clk),
	.d(\internal_counter[22]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[22]~q ),
	.prn(vcc));
defparam \counter_snapshot[22] .is_wysiwyg = "true";
defparam \counter_snapshot[22] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[6]~19 (
	.dataa(\read_mux_out[6]~17_combout ),
	.datab(\read_mux_out~18_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[22]~q ),
	.cin(gnd),
	.combout(\read_mux_out[6]~19_combout ),
	.cout());
defparam \read_mux_out[6]~19 .lut_mask = 16'hFFFE;
defparam \read_mux_out[6]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[7]~20 (
	.dataa(\Equal6~3_combout ),
	.datab(\period_h_register[7]~q ),
	.datac(\Equal6~2_combout ),
	.datad(\period_l_register[7]~q ),
	.cin(gnd),
	.combout(\read_mux_out[7]~20_combout ),
	.cout());
defparam \read_mux_out[7]~20 .lut_mask = 16'hFEFF;
defparam \read_mux_out[7]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter_snapshot[7]~6 (
	.dataa(\internal_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[7]~6_combout ),
	.cout());
defparam \counter_snapshot[7]~6 .lut_mask = 16'h5555;
defparam \counter_snapshot[7]~6 .sum_lutc_input = "datac";

dffeas \counter_snapshot[7] (
	.clk(clk),
	.d(\counter_snapshot[7]~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[7]~q ),
	.prn(vcc));
defparam \counter_snapshot[7] .is_wysiwyg = "true";
defparam \counter_snapshot[7] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~21 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[7]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~21_combout ),
	.cout());
defparam \read_mux_out~21 .lut_mask = 16'hEFFF;
defparam \read_mux_out~21 .sum_lutc_input = "datac";

dffeas \counter_snapshot[23] (
	.clk(clk),
	.d(\internal_counter[23]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[23]~q ),
	.prn(vcc));
defparam \counter_snapshot[23] .is_wysiwyg = "true";
defparam \counter_snapshot[23] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[7]~22 (
	.dataa(\read_mux_out[7]~20_combout ),
	.datab(\read_mux_out~21_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[23]~q ),
	.cin(gnd),
	.combout(\read_mux_out[7]~22_combout ),
	.cout());
defparam \read_mux_out[7]~22 .lut_mask = 16'hFFFE;
defparam \read_mux_out[7]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[15]~23 (
	.dataa(\Equal6~3_combout ),
	.datab(\period_h_register[15]~q ),
	.datac(\Equal6~2_combout ),
	.datad(\period_l_register[15]~q ),
	.cin(gnd),
	.combout(\read_mux_out[15]~23_combout ),
	.cout());
defparam \read_mux_out[15]~23 .lut_mask = 16'hFEFF;
defparam \read_mux_out[15]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter_snapshot[15]~7 (
	.dataa(\internal_counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[15]~7_combout ),
	.cout());
defparam \counter_snapshot[15]~7 .lut_mask = 16'h5555;
defparam \counter_snapshot[15]~7 .sum_lutc_input = "datac";

dffeas \counter_snapshot[15] (
	.clk(clk),
	.d(\counter_snapshot[15]~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[15]~q ),
	.prn(vcc));
defparam \counter_snapshot[15] .is_wysiwyg = "true";
defparam \counter_snapshot[15] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~24 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[15]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~24_combout ),
	.cout());
defparam \read_mux_out~24 .lut_mask = 16'hEFFF;
defparam \read_mux_out~24 .sum_lutc_input = "datac";

dffeas \counter_snapshot[31] (
	.clk(clk),
	.d(\internal_counter[31]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[31]~q ),
	.prn(vcc));
defparam \counter_snapshot[31] .is_wysiwyg = "true";
defparam \counter_snapshot[31] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[15]~25 (
	.dataa(\read_mux_out[15]~23_combout ),
	.datab(\read_mux_out~24_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[31]~q ),
	.cin(gnd),
	.combout(\read_mux_out[15]~25_combout ),
	.cout());
defparam \read_mux_out[15]~25 .lut_mask = 16'hFFFE;
defparam \read_mux_out[15]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[14]~26 (
	.dataa(\Equal6~2_combout ),
	.datab(\Equal6~3_combout ),
	.datac(\period_h_register[14]~q ),
	.datad(\period_l_register[14]~q ),
	.cin(gnd),
	.combout(\read_mux_out[14]~26_combout ),
	.cout());
defparam \read_mux_out[14]~26 .lut_mask = 16'hFFFE;
defparam \read_mux_out[14]~26 .sum_lutc_input = "datac";

dffeas \counter_snapshot[14] (
	.clk(clk),
	.d(\internal_counter[14]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[14]~q ),
	.prn(vcc));
defparam \counter_snapshot[14] .is_wysiwyg = "true";
defparam \counter_snapshot[14] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~27 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[14]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~27_combout ),
	.cout());
defparam \read_mux_out~27 .lut_mask = 16'hEFFF;
defparam \read_mux_out~27 .sum_lutc_input = "datac";

dffeas \counter_snapshot[30] (
	.clk(clk),
	.d(\internal_counter[30]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[30]~q ),
	.prn(vcc));
defparam \counter_snapshot[30] .is_wysiwyg = "true";
defparam \counter_snapshot[30] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[14]~28 (
	.dataa(\read_mux_out[14]~26_combout ),
	.datab(\read_mux_out~27_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[30]~q ),
	.cin(gnd),
	.combout(\read_mux_out[14]~28_combout ),
	.cout());
defparam \read_mux_out[14]~28 .lut_mask = 16'hFFFE;
defparam \read_mux_out[14]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[13]~29 (
	.dataa(\Equal6~2_combout ),
	.datab(\Equal6~3_combout ),
	.datac(\period_h_register[13]~q ),
	.datad(\period_l_register[13]~q ),
	.cin(gnd),
	.combout(\read_mux_out[13]~29_combout ),
	.cout());
defparam \read_mux_out[13]~29 .lut_mask = 16'hFFFE;
defparam \read_mux_out[13]~29 .sum_lutc_input = "datac";

dffeas \counter_snapshot[13] (
	.clk(clk),
	.d(\internal_counter[13]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[13]~q ),
	.prn(vcc));
defparam \counter_snapshot[13] .is_wysiwyg = "true";
defparam \counter_snapshot[13] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~30 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[13]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~30_combout ),
	.cout());
defparam \read_mux_out~30 .lut_mask = 16'hEFFF;
defparam \read_mux_out~30 .sum_lutc_input = "datac";

dffeas \counter_snapshot[29] (
	.clk(clk),
	.d(\internal_counter[29]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[29]~q ),
	.prn(vcc));
defparam \counter_snapshot[29] .is_wysiwyg = "true";
defparam \counter_snapshot[29] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[13]~31 (
	.dataa(\read_mux_out[13]~29_combout ),
	.datab(\read_mux_out~30_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[29]~q ),
	.cin(gnd),
	.combout(\read_mux_out[13]~31_combout ),
	.cout());
defparam \read_mux_out[13]~31 .lut_mask = 16'hFFFE;
defparam \read_mux_out[13]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[12]~32 (
	.dataa(\Equal6~2_combout ),
	.datab(\Equal6~3_combout ),
	.datac(\period_h_register[12]~q ),
	.datad(\period_l_register[12]~q ),
	.cin(gnd),
	.combout(\read_mux_out[12]~32_combout ),
	.cout());
defparam \read_mux_out[12]~32 .lut_mask = 16'hFFFE;
defparam \read_mux_out[12]~32 .sum_lutc_input = "datac";

dffeas \counter_snapshot[12] (
	.clk(clk),
	.d(\internal_counter[12]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[12]~q ),
	.prn(vcc));
defparam \counter_snapshot[12] .is_wysiwyg = "true";
defparam \counter_snapshot[12] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~33 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[12]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~33_combout ),
	.cout());
defparam \read_mux_out~33 .lut_mask = 16'hEFFF;
defparam \read_mux_out~33 .sum_lutc_input = "datac";

dffeas \counter_snapshot[28] (
	.clk(clk),
	.d(\internal_counter[28]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[28]~q ),
	.prn(vcc));
defparam \counter_snapshot[28] .is_wysiwyg = "true";
defparam \counter_snapshot[28] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[12]~34 (
	.dataa(\read_mux_out[12]~32_combout ),
	.datab(\read_mux_out~33_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[28]~q ),
	.cin(gnd),
	.combout(\read_mux_out[12]~34_combout ),
	.cout());
defparam \read_mux_out[12]~34 .lut_mask = 16'hFFFE;
defparam \read_mux_out[12]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[11]~35 (
	.dataa(\Equal6~2_combout ),
	.datab(\Equal6~3_combout ),
	.datac(\period_h_register[11]~q ),
	.datad(\period_l_register[11]~q ),
	.cin(gnd),
	.combout(\read_mux_out[11]~35_combout ),
	.cout());
defparam \read_mux_out[11]~35 .lut_mask = 16'hFFFE;
defparam \read_mux_out[11]~35 .sum_lutc_input = "datac";

dffeas \counter_snapshot[11] (
	.clk(clk),
	.d(\internal_counter[11]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[11]~q ),
	.prn(vcc));
defparam \counter_snapshot[11] .is_wysiwyg = "true";
defparam \counter_snapshot[11] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~36 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[11]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~36_combout ),
	.cout());
defparam \read_mux_out~36 .lut_mask = 16'hEFFF;
defparam \read_mux_out~36 .sum_lutc_input = "datac";

dffeas \counter_snapshot[27] (
	.clk(clk),
	.d(\internal_counter[27]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[27]~q ),
	.prn(vcc));
defparam \counter_snapshot[27] .is_wysiwyg = "true";
defparam \counter_snapshot[27] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[11]~37 (
	.dataa(\read_mux_out[11]~35_combout ),
	.datab(\read_mux_out~36_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[27]~q ),
	.cin(gnd),
	.combout(\read_mux_out[11]~37_combout ),
	.cout());
defparam \read_mux_out[11]~37 .lut_mask = 16'hFFFE;
defparam \read_mux_out[11]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[10]~38 (
	.dataa(\Equal6~3_combout ),
	.datab(\period_h_register[10]~q ),
	.datac(\Equal6~2_combout ),
	.datad(\period_l_register[10]~q ),
	.cin(gnd),
	.combout(\read_mux_out[10]~38_combout ),
	.cout());
defparam \read_mux_out[10]~38 .lut_mask = 16'hFEFF;
defparam \read_mux_out[10]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter_snapshot[10]~8 (
	.dataa(\internal_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[10]~8_combout ),
	.cout());
defparam \counter_snapshot[10]~8 .lut_mask = 16'h5555;
defparam \counter_snapshot[10]~8 .sum_lutc_input = "datac";

dffeas \counter_snapshot[10] (
	.clk(clk),
	.d(\counter_snapshot[10]~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[10]~q ),
	.prn(vcc));
defparam \counter_snapshot[10] .is_wysiwyg = "true";
defparam \counter_snapshot[10] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~39 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[10]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~39_combout ),
	.cout());
defparam \read_mux_out~39 .lut_mask = 16'hEFFF;
defparam \read_mux_out~39 .sum_lutc_input = "datac";

dffeas \counter_snapshot[26] (
	.clk(clk),
	.d(\internal_counter[26]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[26]~q ),
	.prn(vcc));
defparam \counter_snapshot[26] .is_wysiwyg = "true";
defparam \counter_snapshot[26] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[10]~40 (
	.dataa(\read_mux_out[10]~38_combout ),
	.datab(\read_mux_out~39_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[26]~q ),
	.cin(gnd),
	.combout(\read_mux_out[10]~40_combout ),
	.cout());
defparam \read_mux_out[10]~40 .lut_mask = 16'hFFFE;
defparam \read_mux_out[10]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[9]~41 (
	.dataa(\Equal6~3_combout ),
	.datab(\period_h_register[9]~q ),
	.datac(\Equal6~2_combout ),
	.datad(\period_l_register[9]~q ),
	.cin(gnd),
	.combout(\read_mux_out[9]~41_combout ),
	.cout());
defparam \read_mux_out[9]~41 .lut_mask = 16'hFEFF;
defparam \read_mux_out[9]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter_snapshot[9]~9 (
	.dataa(\internal_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter_snapshot[9]~9_combout ),
	.cout());
defparam \counter_snapshot[9]~9 .lut_mask = 16'h5555;
defparam \counter_snapshot[9]~9 .sum_lutc_input = "datac";

dffeas \counter_snapshot[9] (
	.clk(clk),
	.d(\counter_snapshot[9]~9_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[9]~q ),
	.prn(vcc));
defparam \counter_snapshot[9] .is_wysiwyg = "true";
defparam \counter_snapshot[9] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~42 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[9]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~42_combout ),
	.cout());
defparam \read_mux_out~42 .lut_mask = 16'hEFFF;
defparam \read_mux_out~42 .sum_lutc_input = "datac";

dffeas \counter_snapshot[25] (
	.clk(clk),
	.d(\internal_counter[25]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[25]~q ),
	.prn(vcc));
defparam \counter_snapshot[25] .is_wysiwyg = "true";
defparam \counter_snapshot[25] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[9]~43 (
	.dataa(\read_mux_out[9]~41_combout ),
	.datab(\read_mux_out~42_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[25]~q ),
	.cin(gnd),
	.combout(\read_mux_out[9]~43_combout ),
	.cout());
defparam \read_mux_out[9]~43 .lut_mask = 16'hFFFE;
defparam \read_mux_out[9]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[8]~44 (
	.dataa(\Equal6~2_combout ),
	.datab(\Equal6~3_combout ),
	.datac(\period_h_register[8]~q ),
	.datad(\period_l_register[8]~q ),
	.cin(gnd),
	.combout(\read_mux_out[8]~44_combout ),
	.cout());
defparam \read_mux_out[8]~44 .lut_mask = 16'hFFFE;
defparam \read_mux_out[8]~44 .sum_lutc_input = "datac";

dffeas \counter_snapshot[8] (
	.clk(clk),
	.d(\internal_counter[8]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[8]~q ),
	.prn(vcc));
defparam \counter_snapshot[8] .is_wysiwyg = "true";
defparam \counter_snapshot[8] .power_up = "low";

cycloneive_lcell_comb \read_mux_out~45 (
	.dataa(W_alu_result_4),
	.datab(\counter_snapshot[8]~q ),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\read_mux_out~45_combout ),
	.cout());
defparam \read_mux_out~45 .lut_mask = 16'hEFFF;
defparam \read_mux_out~45 .sum_lutc_input = "datac";

dffeas \counter_snapshot[24] (
	.clk(clk),
	.d(\internal_counter[24]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[24]~q ),
	.prn(vcc));
defparam \counter_snapshot[24] .is_wysiwyg = "true";
defparam \counter_snapshot[24] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[8]~46 (
	.dataa(\read_mux_out[8]~44_combout ),
	.datab(\read_mux_out~45_combout ),
	.datac(\Equal6~4_combout ),
	.datad(\counter_snapshot[24]~q ),
	.cin(gnd),
	.combout(\read_mux_out[8]~46_combout ),
	.cout());
defparam \read_mux_out[8]~46 .lut_mask = 16'hFFFE;
defparam \read_mux_out[8]~46 .sum_lutc_input = "datac";

endmodule
